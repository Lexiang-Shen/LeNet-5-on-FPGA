`define LINEAR2_WEIGHT \
reg [0:17] linear2_weight_array [0:9][0:11];\
always@(posedge clk) begin\
    linear2_weight_array[0][0] <= 18'h000c9;\
    linear2_weight_array[0][1] <= 18'h200b1;\
    linear2_weight_array[0][2] <= 18'h200b7;\
    linear2_weight_array[0][3] <= 18'h001d3;\
    linear2_weight_array[0][4] <= 18'h200d5;\
    linear2_weight_array[0][5] <= 18'h202a7;\
    linear2_weight_array[0][6] <= 18'h2019f;\
    linear2_weight_array[0][7] <= 18'h2009a;\
    linear2_weight_array[0][8] <= 18'h20096;\
    linear2_weight_array[0][9] <= 18'h000da;\
    linear2_weight_array[0][10] <= 18'h2010d;\
    linear2_weight_array[0][11] <= 18'h0008c;\
    linear2_weight_array[1][0] <= 18'h20315;\
    linear2_weight_array[1][1] <= 18'h20087;\
    linear2_weight_array[1][2] <= 18'h001cb;\
    linear2_weight_array[1][3] <= 18'h20246;\
    linear2_weight_array[1][4] <= 18'h000c6;\
    linear2_weight_array[1][5] <= 18'h0001d;\
    linear2_weight_array[1][6] <= 18'h00080;\
    linear2_weight_array[1][7] <= 18'h20112;\
    linear2_weight_array[1][8] <= 18'h200a5;\
    linear2_weight_array[1][9] <= 18'h0016f;\
    linear2_weight_array[1][10] <= 18'h200b0;\
    linear2_weight_array[1][11] <= 18'h000c5;\
    linear2_weight_array[2][0] <= 18'h00069;\
    linear2_weight_array[2][1] <= 18'h2009d;\
    linear2_weight_array[2][2] <= 18'h0019e;\
    linear2_weight_array[2][3] <= 18'h20221;\
    linear2_weight_array[2][4] <= 18'h20071;\
    linear2_weight_array[2][5] <= 18'h2022b;\
    linear2_weight_array[2][6] <= 18'h20155;\
    linear2_weight_array[2][7] <= 18'h000c1;\
    linear2_weight_array[2][8] <= 18'h200d1;\
    linear2_weight_array[2][9] <= 18'h201d0;\
    linear2_weight_array[2][10] <= 18'h000c5;\
    linear2_weight_array[2][11] <= 18'h00132;\
    linear2_weight_array[3][0] <= 18'h000bb;\
    linear2_weight_array[3][1] <= 18'h200ad;\
    linear2_weight_array[3][2] <= 18'h00047;\
    linear2_weight_array[3][3] <= 18'h20237;\
    linear2_weight_array[3][4] <= 18'h200e8;\
    linear2_weight_array[3][5] <= 18'h000a4;\
    linear2_weight_array[3][6] <= 18'h200dc;\
    linear2_weight_array[3][7] <= 18'h20127;\
    linear2_weight_array[3][8] <= 18'h00007;\
    linear2_weight_array[3][9] <= 18'h0004c;\
    linear2_weight_array[3][10] <= 18'h00010;\
    linear2_weight_array[3][11] <= 18'h00121;\
    linear2_weight_array[4][0] <= 18'h201fd;\
    linear2_weight_array[4][1] <= 18'h000f5;\
    linear2_weight_array[4][2] <= 18'h2017b;\
    linear2_weight_array[4][3] <= 18'h00022;\
    linear2_weight_array[4][4] <= 18'h00006;\
    linear2_weight_array[4][5] <= 18'h001f5;\
    linear2_weight_array[4][6] <= 18'h2001a;\
    linear2_weight_array[4][7] <= 18'h0023f;\
    linear2_weight_array[4][8] <= 18'h000ed;\
    linear2_weight_array[4][9] <= 18'h201a7;\
    linear2_weight_array[4][10] <= 18'h20064;\
    linear2_weight_array[4][11] <= 18'h0009e;\
    linear2_weight_array[5][0] <= 18'h00171;\
    linear2_weight_array[5][1] <= 18'h000b6;\
    linear2_weight_array[5][2] <= 18'h20095;\
    linear2_weight_array[5][3] <= 18'h200ed;\
    linear2_weight_array[5][4] <= 18'h00026;\
    linear2_weight_array[5][5] <= 18'h00188;\
    linear2_weight_array[5][6] <= 18'h201ac;\
    linear2_weight_array[5][7] <= 18'h201c8;\
    linear2_weight_array[5][8] <= 18'h00024;\
    linear2_weight_array[5][9] <= 18'h200e5;\
    linear2_weight_array[5][10] <= 18'h00005;\
    linear2_weight_array[5][11] <= 18'h20169;\
    linear2_weight_array[6][0] <= 18'h0003d;\
    linear2_weight_array[6][1] <= 18'h2000b;\
    linear2_weight_array[6][2] <= 18'h00081;\
    linear2_weight_array[6][3] <= 18'h0019a;\
    linear2_weight_array[6][4] <= 18'h200ed;\
    linear2_weight_array[6][5] <= 18'h0008a;\
    linear2_weight_array[6][6] <= 18'h202c5;\
    linear2_weight_array[6][7] <= 18'h0000b;\
    linear2_weight_array[6][8] <= 18'h2006d;\
    linear2_weight_array[6][9] <= 18'h20068;\
    linear2_weight_array[6][10] <= 18'h20082;\
    linear2_weight_array[6][11] <= 18'h20308;\
    linear2_weight_array[7][0] <= 18'h0001e;\
    linear2_weight_array[7][1] <= 18'h2007f;\
    linear2_weight_array[7][2] <= 18'h0002e;\
    linear2_weight_array[7][3] <= 18'h20110;\
    linear2_weight_array[7][4] <= 18'h2006c;\
    linear2_weight_array[7][5] <= 18'h20104;\
    linear2_weight_array[7][6] <= 18'h00234;\
    linear2_weight_array[7][7] <= 18'h2003a;\
    linear2_weight_array[7][8] <= 18'h20081;\
    linear2_weight_array[7][9] <= 18'h20238;\
    linear2_weight_array[7][10] <= 18'h20054;\
    linear2_weight_array[7][11] <= 18'h20047;\
    linear2_weight_array[8][0] <= 18'h000df;\
    linear2_weight_array[8][1] <= 18'h000f6;\
    linear2_weight_array[8][2] <= 18'h20005;\
    linear2_weight_array[8][3] <= 18'h20158;\
    linear2_weight_array[8][4] <= 18'h0001c;\
    linear2_weight_array[8][5] <= 18'h200a2;\
    linear2_weight_array[8][6] <= 18'h20177;\
    linear2_weight_array[8][7] <= 18'h0015b;\
    linear2_weight_array[8][8] <= 18'h0010c;\
    linear2_weight_array[8][9] <= 18'h00143;\
    linear2_weight_array[8][10] <= 18'h00081;\
    linear2_weight_array[8][11] <= 18'h201b0;\
    linear2_weight_array[9][0] <= 18'h00065;\
    linear2_weight_array[9][1] <= 18'h200ce;\
    linear2_weight_array[9][2] <= 18'h20366;\
    linear2_weight_array[9][3] <= 18'h2006f;\
    linear2_weight_array[9][4] <= 18'h200d4;\
    linear2_weight_array[9][5] <= 18'h00011;\
    linear2_weight_array[9][6] <= 18'h00097;\
    linear2_weight_array[9][7] <= 18'h00159;\
    linear2_weight_array[9][8] <= 18'h200b9;\
    linear2_weight_array[9][9] <= 18'h00041;\
    linear2_weight_array[9][10] <= 18'h00030;\
    linear2_weight_array[9][11] <= 18'h00090;\
end

/*
`define LINEAR2_WEIGHT \
reg [0:18] linear2_weight_array [0:9][0:11];\
always@(posedge clk or negedge rst_n) begin\
    linear2_weight_array[0][ 0] <= 18'h01000;\
    linear2_weight_array[0][ 1] <= 18'h20300;\
    linear2_weight_array[0][ 2] <= 18'h00d00;\
    linear2_weight_array[0][ 3] <= 18'h22800;\
    linear2_weight_array[0][ 4] <= 18'h01000;\
    linear2_weight_array[0][ 5] <= 18'h20300;\
    linear2_weight_array[0][ 6] <= 18'h00d00;\
    linear2_weight_array[0][ 7] <= 18'h22800;\
    linear2_weight_array[0][ 8] <= 18'h01000;\
    linear2_weight_array[0][ 9] <= 18'h20300;\
    linear2_weight_array[0][10] <= 18'h00d00;\
    linear2_weight_array[0][11] <= 18'h22800;\
    linear2_weight_array[1][ 0] <= 18'h00c00;\
    linear2_weight_array[1][ 1] <= 18'h00500;\
    linear2_weight_array[1][ 2] <= 18'h21300;\
    linear2_weight_array[1][ 3] <= 18'h00280;\
    linear2_weight_array[1][ 4] <= 18'h00c00;\
    linear2_weight_array[1][ 5] <= 18'h00500;\
    linear2_weight_array[1][ 6] <= 18'h21300;\
    linear2_weight_array[1][ 7] <= 18'h00280;\
    linear2_weight_array[1][ 8] <= 18'h00c00;\
    linear2_weight_array[1][ 9] <= 18'h00500;\
    linear2_weight_array[1][10] <= 18'h21300;\
    linear2_weight_array[1][11] <= 18'h00280;\
    linear2_weight_array[2][ 0] <= 18'h01000;\
    linear2_weight_array[2][ 1] <= 18'h20300;\
    linear2_weight_array[2][ 2] <= 18'h00d00;\
    linear2_weight_array[2][ 3] <= 18'h22800;\
    linear2_weight_array[2][ 4] <= 18'h01000;\
    linear2_weight_array[2][ 5] <= 18'h20300;\
    linear2_weight_array[2][ 6] <= 18'h00d00;\
    linear2_weight_array[2][ 7] <= 18'h22800;\
    linear2_weight_array[2][ 8] <= 18'h01000;\
    linear2_weight_array[2][ 9] <= 18'h20300;\
    linear2_weight_array[2][10] <= 18'h00d00;\
    linear2_weight_array[2][11] <= 18'h22800;\
    linear2_weight_array[3][ 0] <= 18'h00c00;\
    linear2_weight_array[3][ 1] <= 18'h00500;\
    linear2_weight_array[3][ 2] <= 18'h21300;\
    linear2_weight_array[3][ 3] <= 18'h00280;\
    linear2_weight_array[3][ 4] <= 18'h00c00;\
    linear2_weight_array[3][ 5] <= 18'h00500;\
    linear2_weight_array[3][ 6] <= 18'h21300;\
    linear2_weight_array[3][ 7] <= 18'h00280;\
    linear2_weight_array[3][ 8] <= 18'h00c00;\
    linear2_weight_array[3][ 9] <= 18'h00500;\
    linear2_weight_array[3][10] <= 18'h21300;\
    linear2_weight_array[3][11] <= 18'h00280;\
    linear2_weight_array[4][ 0] <= 18'h01000;\
    linear2_weight_array[4][ 1] <= 18'h20300;\
    linear2_weight_array[4][ 2] <= 18'h00d00;\
    linear2_weight_array[4][ 3] <= 18'h22800;\
    linear2_weight_array[4][ 4] <= 18'h01000;\
    linear2_weight_array[4][ 5] <= 18'h20300;\
    linear2_weight_array[4][ 6] <= 18'h00d00;\
    linear2_weight_array[4][ 7] <= 18'h22800;\
    linear2_weight_array[4][ 8] <= 18'h01000;\
    linear2_weight_array[4][ 9] <= 18'h20300;\
    linear2_weight_array[4][10] <= 18'h00d00;\
    linear2_weight_array[4][11] <= 18'h22800;\
    linear2_weight_array[5][ 0] <= 18'h00c00;\
    linear2_weight_array[5][ 1] <= 18'h00500;\
    linear2_weight_array[5][ 2] <= 18'h21300;\
    linear2_weight_array[5][ 3] <= 18'h00280;\
    linear2_weight_array[5][ 4] <= 18'h00c00;\
    linear2_weight_array[5][ 5] <= 18'h00500;\
    linear2_weight_array[5][ 6] <= 18'h21300;\
    linear2_weight_array[5][ 7] <= 18'h00280;\
    linear2_weight_array[5][ 8] <= 18'h00c00;\
    linear2_weight_array[5][ 9] <= 18'h00500;\
    linear2_weight_array[5][10] <= 18'h21300;\
    linear2_weight_array[5][11] <= 18'h00280;\
    linear2_weight_array[6][ 0] <= 18'h01000;\
    linear2_weight_array[6][ 1] <= 18'h20300;\
    linear2_weight_array[6][ 2] <= 18'h00d00;\
    linear2_weight_array[6][ 3] <= 18'h22800;\
    linear2_weight_array[6][ 4] <= 18'h01000;\
    linear2_weight_array[6][ 5] <= 18'h20300;\
    linear2_weight_array[6][ 6] <= 18'h00d00;\
    linear2_weight_array[6][ 7] <= 18'h22800;\
    linear2_weight_array[6][ 8] <= 18'h01000;\
    linear2_weight_array[6][ 9] <= 18'h20300;\
    linear2_weight_array[6][10] <= 18'h00d00;\
    linear2_weight_array[6][11] <= 18'h22800;\
    linear2_weight_array[7][ 0] <= 18'h00c00;\
    linear2_weight_array[7][ 1] <= 18'h00500;\
    linear2_weight_array[7][ 2] <= 18'h21300;\
    linear2_weight_array[7][ 3] <= 18'h00280;\
    linear2_weight_array[7][ 4] <= 18'h00c00;\
    linear2_weight_array[7][ 5] <= 18'h00500;\
    linear2_weight_array[7][ 6] <= 18'h21300;\
    linear2_weight_array[7][ 7] <= 18'h00280;\
    linear2_weight_array[7][ 8] <= 18'h00c00;\
    linear2_weight_array[7][ 9] <= 18'h00500;\
    linear2_weight_array[7][10] <= 18'h21300;\
    linear2_weight_array[7][11] <= 18'h00280;\
    linear2_weight_array[8][ 0] <= 18'h01000;\
    linear2_weight_array[8][ 1] <= 18'h20300;\
    linear2_weight_array[8][ 2] <= 18'h00d00;\
    linear2_weight_array[8][ 3] <= 18'h22800;\
    linear2_weight_array[8][ 4] <= 18'h01000;\
    linear2_weight_array[8][ 5] <= 18'h20300;\
    linear2_weight_array[8][ 6] <= 18'h00d00;\
    linear2_weight_array[8][ 7] <= 18'h22800;\
    linear2_weight_array[8][ 8] <= 18'h01000;\
    linear2_weight_array[8][ 9] <= 18'h20300;\
    linear2_weight_array[8][10] <= 18'h00d00;\
    linear2_weight_array[8][11] <= 18'h22800;\
    linear2_weight_array[9][ 0] <= 18'h00c00;\
    linear2_weight_array[9][ 1] <= 18'h00500;\
    linear2_weight_array[9][ 2] <= 18'h21300;\
    linear2_weight_array[9][ 3] <= 18'h00280;\
    linear2_weight_array[9][ 4] <= 18'h00c00;\
    linear2_weight_array[9][ 5] <= 18'h00500;\
    linear2_weight_array[9][ 6] <= 18'h21300;\
    linear2_weight_array[9][ 7] <= 18'h00280;\
    linear2_weight_array[9][ 8] <= 18'h00c00;\
    linear2_weight_array[9][ 9] <= 18'h00500;\
    linear2_weight_array[9][10] <= 18'h21300;\
    linear2_weight_array[9][11] <= 18'h00280;\
end
*/