`define ADDED \
always@(posedge clk or negedge rst_n) begin\
    if(!rst_n) begin\
		added_1[0] <= 18'd0;\
		added_1[1] <= 18'd0;\
		added_1[2] <= 18'd0;\
		added_1[3] <= 18'd0;\
		added_1[4] <= 18'd0;\
		added_1[5] <= 18'd0;\
		added_1[6] <= 18'd0;\
		added_1[7] <= 18'd0;\
		added_1[8] <= 18'd0;\
		added_1[9] <= 18'd0;\
		added_1[10] <= 18'd0;\
		added_1[11] <= 18'd0;\
		added_1[12] <= 18'd0;\
		added_1[13] <= 18'd0;\
		added_1[14] <= 18'd0;\
		added_1[15] <= 18'd0;\
		added_1[16] <= 18'd0;\
		added_1[17] <= 18'd0;\
		added_1[18] <= 18'd0;\
		added_1[19] <= 18'd0;\
		added_1[20] <= 18'd0;\
		added_1[21] <= 18'd0;\
		added_1[22] <= 18'd0;\
		added_1[23] <= 18'd0;\
		added_1[24] <= 18'd0;\
		added_1[25] <= 18'd0;\
		added_1[26] <= 18'd0;\
		added_1[27] <= 18'd0;\
		added_1[28] <= 18'd0;\
		added_1[29] <= 18'd0;\
		added_1[30] <= 18'd0;\
		added_1[31] <= 18'd0;\
		added_1[32] <= 18'd0;\
		added_1[33] <= 18'd0;\
		added_1[34] <= 18'd0;\
		added_1[35] <= 18'd0;\
		added_1[36] <= 18'd0;\
		added_1[37] <= 18'd0;\
		added_1[38] <= 18'd0;\
		added_1[39] <= 18'd0;\
		added_1[40] <= 18'd0;\
		added_1[41] <= 18'd0;\
		added_1[42] <= 18'd0;\
		added_1[43] <= 18'd0;\
		added_1[44] <= 18'd0;\
		added_1[45] <= 18'd0;\
		added_1[46] <= 18'd0;\
		added_1[47] <= 18'd0;\
		added_1[48] <= 18'd0;\
		added_1[49] <= 18'd0;\
		added_1[50] <= 18'd0;\
		added_1[51] <= 18'd0;\
		added_1[52] <= 18'd0;\
		added_1[53] <= 18'd0;\
		added_1[54] <= 18'd0;\
		added_1[55] <= 18'd0;\
		added_1[56] <= 18'd0;\
		added_1[57] <= 18'd0;\
		added_1[58] <= 18'd0;\
		added_1[59] <= 18'd0;\
		added_1[60] <= 18'd0;\
		added_1[61] <= 18'd0;\
		added_1[62] <= 18'd0;\
		added_1[63] <= 18'd0;\
		added_1[64] <= 18'd0;\
		added_1[65] <= 18'd0;\
		added_1[66] <= 18'd0;\
		added_1[67] <= 18'd0;\
		added_1[68] <= 18'd0;\
		added_1[69] <= 18'd0;\
		added_1[70] <= 18'd0;\
		added_1[71] <= 18'd0;\
		added_1[72] <= 18'd0;\
		added_1[73] <= 18'd0;\
		added_1[74] <= 18'd0;\
		added_1[75] <= 18'd0;\
		added_1[76] <= 18'd0;\
		added_1[77] <= 18'd0;\
		added_1[78] <= 18'd0;\
		added_1[79] <= 18'd0;\
		added_1[80] <= 18'd0;\
		added_1[81] <= 18'd0;\
		added_1[82] <= 18'd0;\
		added_1[83] <= 18'd0;\
		added_1[84] <= 18'd0;\
		added_1[85] <= 18'd0;\
		added_1[86] <= 18'd0;\
		added_1[87] <= 18'd0;\
		added_1[88] <= 18'd0;\
		added_1[89] <= 18'd0;\
		added_1[90] <= 18'd0;\
		added_1[91] <= 18'd0;\
		added_1[92] <= 18'd0;\
		added_1[93] <= 18'd0;\
		added_1[94] <= 18'd0;\
		added_1[95] <= 18'd0;\
		added_1[96] <= 18'd0;\
		added_1[97] <= 18'd0;\
		added_1[98] <= 18'd0;\
		added_1[99] <= 18'd0;\
		added_1[100] <= 18'd0;\
		added_1[101] <= 18'd0;\
		added_1[102] <= 18'd0;\
		added_1[103] <= 18'd0;\
		added_1[104] <= 18'd0;\
		added_1[105] <= 18'd0;\
		added_1[106] <= 18'd0;\
		added_1[107] <= 18'd0;\
		added_1[108] <= 18'd0;\
		added_1[109] <= 18'd0;\
		added_1[110] <= 18'd0;\
		added_1[111] <= 18'd0;\
		added_2[0] <= 18'd0;\
		added_2[1] <= 18'd0;\
		added_2[2] <= 18'd0;\
		added_2[3] <= 18'd0;\
		added_2[4] <= 18'd0;\
		added_2[5] <= 18'd0;\
		added_2[6] <= 18'd0;\
		added_2[7] <= 18'd0;\
		added_2[8] <= 18'd0;\
		added_2[9] <= 18'd0;\
		added_2[10] <= 18'd0;\
		added_2[11] <= 18'd0;\
		added_2[12] <= 18'd0;\
		added_2[13] <= 18'd0;\
		added_2[14] <= 18'd0;\
		added_2[15] <= 18'd0;\
		added_2[16] <= 18'd0;\
		added_2[17] <= 18'd0;\
		added_2[18] <= 18'd0;\
		added_2[19] <= 18'd0;\
		added_2[20] <= 18'd0;\
		added_2[21] <= 18'd0;\
		added_2[22] <= 18'd0;\
		added_2[23] <= 18'd0;\
		added_2[24] <= 18'd0;\
		added_2[25] <= 18'd0;\
		added_2[26] <= 18'd0;\
		added_2[27] <= 18'd0;\
		added_2[28] <= 18'd0;\
		added_2[29] <= 18'd0;\
		added_2[30] <= 18'd0;\
		added_2[31] <= 18'd0;\
		added_2[32] <= 18'd0;\
		added_2[33] <= 18'd0;\
		added_2[34] <= 18'd0;\
		added_2[35] <= 18'd0;\
		added_2[36] <= 18'd0;\
		added_2[37] <= 18'd0;\
		added_2[38] <= 18'd0;\
		added_2[39] <= 18'd0;\
		added_2[40] <= 18'd0;\
		added_2[41] <= 18'd0;\
		added_2[42] <= 18'd0;\
		added_2[43] <= 18'd0;\
		added_2[44] <= 18'd0;\
		added_2[45] <= 18'd0;\
		added_2[46] <= 18'd0;\
		added_2[47] <= 18'd0;\
		added_2[48] <= 18'd0;\
		added_2[49] <= 18'd0;\
		added_2[50] <= 18'd0;\
		added_2[51] <= 18'd0;\
		added_2[52] <= 18'd0;\
		added_2[53] <= 18'd0;\
		added_2[54] <= 18'd0;\
		added_2[55] <= 18'd0;\
		added_2[56] <= 18'd0;\
		added_2[57] <= 18'd0;\
		added_2[58] <= 18'd0;\
		added_2[59] <= 18'd0;\
		added_2[60] <= 18'd0;\
		added_2[61] <= 18'd0;\
		added_2[62] <= 18'd0;\
		added_2[63] <= 18'd0;\
		added_2[64] <= 18'd0;\
		added_2[65] <= 18'd0;\
		added_2[66] <= 18'd0;\
		added_2[67] <= 18'd0;\
		added_2[68] <= 18'd0;\
		added_2[69] <= 18'd0;\
		added_2[70] <= 18'd0;\
		added_2[71] <= 18'd0;\
		added_2[72] <= 18'd0;\
		added_2[73] <= 18'd0;\
		added_2[74] <= 18'd0;\
		added_2[75] <= 18'd0;\
		added_2[76] <= 18'd0;\
		added_2[77] <= 18'd0;\
		added_2[78] <= 18'd0;\
		added_2[79] <= 18'd0;\
		added_2[80] <= 18'd0;\
		added_2[81] <= 18'd0;\
		added_2[82] <= 18'd0;\
		added_2[83] <= 18'd0;\
		added_2[84] <= 18'd0;\
		added_2[85] <= 18'd0;\
		added_2[86] <= 18'd0;\
		added_2[87] <= 18'd0;\
		added_2[88] <= 18'd0;\
		added_2[89] <= 18'd0;\
		added_2[90] <= 18'd0;\
		added_2[91] <= 18'd0;\
		added_2[92] <= 18'd0;\
		added_2[93] <= 18'd0;\
		added_2[94] <= 18'd0;\
		added_2[95] <= 18'd0;\
		added_2[96] <= 18'd0;\
		added_2[97] <= 18'd0;\
		added_2[98] <= 18'd0;\
		added_2[99] <= 18'd0;\
		added_2[100] <= 18'd0;\
		added_2[101] <= 18'd0;\
		added_2[102] <= 18'd0;\
		added_2[103] <= 18'd0;\
		added_2[104] <= 18'd0;\
		added_2[105] <= 18'd0;\
		added_2[106] <= 18'd0;\
		added_2[107] <= 18'd0;\
		added_2[108] <= 18'd0;\
		added_2[109] <= 18'd0;\
		added_2[110] <= 18'd0;\
		added_2[111] <= 18'd0;\
    end\
    else begin\
        case(state)\
            IDLE     :;\
            INPUT    :;\
            CONV1_1_1,CONV1_1_2,CONV1_1_3,CONV1_1_4,CONV1_1_5,CONV1_1_6,CONV1_1_7:begin \
                if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[0] <= conv1_bias_array[0];\
					added_1[1] <= conv1_bias_array[0];\
					added_1[2] <= conv1_bias_array[0];\
					added_1[3] <= conv1_bias_array[0];\
					added_1[4] <= conv1_bias_array[0];\
					added_1[5] <= conv1_bias_array[0];\
					added_1[6] <= conv1_bias_array[0];\
					added_1[7] <= conv1_bias_array[0];\
					added_1[8] <= conv1_bias_array[0];\
					added_1[9] <= conv1_bias_array[0];\
					added_1[10] <= conv1_bias_array[0];\
					added_1[11] <= conv1_bias_array[0];\
					added_1[12] <= conv1_bias_array[0];\
					added_1[13] <= conv1_bias_array[0];\
					added_1[14] <= conv1_bias_array[0];\
					added_1[15] <= conv1_bias_array[0];\
					added_1[16] <= conv1_bias_array[0];\
					added_1[17] <= conv1_bias_array[0];\
					added_1[18] <= conv1_bias_array[0];\
					added_1[19] <= conv1_bias_array[0];\
					added_1[20] <= conv1_bias_array[0];\
					added_1[21] <= conv1_bias_array[0];\
					added_1[22] <= conv1_bias_array[0];\
					added_1[23] <= conv1_bias_array[0];\
					added_1[24] <= conv1_bias_array[0];\
					added_1[25] <= conv1_bias_array[0];\
					added_1[26] <= conv1_bias_array[0];\
					added_1[27] <= conv1_bias_array[0];\
					added_1[28] <= conv1_bias_array[0];\
					added_1[29] <= conv1_bias_array[0];\
					added_1[30] <= conv1_bias_array[0];\
					added_1[31] <= conv1_bias_array[0];\
					added_1[32] <= conv1_bias_array[0];\
					added_1[33] <= conv1_bias_array[0];\
					added_1[34] <= conv1_bias_array[0];\
					added_1[35] <= conv1_bias_array[0];\
					added_1[36] <= conv1_bias_array[0];\
					added_1[37] <= conv1_bias_array[0];\
					added_1[38] <= conv1_bias_array[0];\
					added_1[39] <= conv1_bias_array[0];\
					added_1[40] <= conv1_bias_array[0];\
					added_1[41] <= conv1_bias_array[0];\
					added_1[42] <= conv1_bias_array[0];\
					added_1[43] <= conv1_bias_array[0];\
					added_1[44] <= conv1_bias_array[0];\
					added_1[45] <= conv1_bias_array[0];\
					added_1[46] <= conv1_bias_array[0];\
					added_1[47] <= conv1_bias_array[0];\
					added_1[48] <= conv1_bias_array[0];\
					added_1[49] <= conv1_bias_array[0];\
					added_1[50] <= conv1_bias_array[0];\
					added_1[51] <= conv1_bias_array[0];\
					added_1[52] <= conv1_bias_array[0];\
					added_1[53] <= conv1_bias_array[0];\
					added_1[54] <= conv1_bias_array[0];\
					added_1[55] <= conv1_bias_array[0];\
					added_1[56] <= conv1_bias_array[0];\
					added_1[57] <= conv1_bias_array[0];\
					added_1[58] <= conv1_bias_array[0];\
					added_1[59] <= conv1_bias_array[0];\
					added_1[60] <= conv1_bias_array[0];\
					added_1[61] <= conv1_bias_array[0];\
					added_1[62] <= conv1_bias_array[0];\
					added_1[63] <= conv1_bias_array[0];\
					added_1[64] <= conv1_bias_array[0];\
					added_1[65] <= conv1_bias_array[0];\
					added_1[66] <= conv1_bias_array[0];\
					added_1[67] <= conv1_bias_array[0];\
					added_1[68] <= conv1_bias_array[0];\
					added_1[69] <= conv1_bias_array[0];\
					added_1[70] <= conv1_bias_array[0];\
					added_1[71] <= conv1_bias_array[0];\
					added_1[72] <= conv1_bias_array[0];\
					added_1[73] <= conv1_bias_array[0];\
					added_1[74] <= conv1_bias_array[0];\
					added_1[75] <= conv1_bias_array[0];\
					added_1[76] <= conv1_bias_array[0];\
					added_1[77] <= conv1_bias_array[0];\
					added_1[78] <= conv1_bias_array[0];\
					added_1[79] <= conv1_bias_array[0];\
					added_1[80] <= conv1_bias_array[0];\
					added_1[81] <= conv1_bias_array[0];\
					added_1[82] <= conv1_bias_array[0];\
					added_1[83] <= conv1_bias_array[0];\
					added_1[84] <= conv1_bias_array[0];\
					added_1[85] <= conv1_bias_array[0];\
					added_1[86] <= conv1_bias_array[0];\
					added_1[87] <= conv1_bias_array[0];\
					added_1[88] <= conv1_bias_array[0];\
					added_1[89] <= conv1_bias_array[0];\
					added_1[90] <= conv1_bias_array[0];\
					added_1[91] <= conv1_bias_array[0];\
					added_1[92] <= conv1_bias_array[0];\
					added_1[93] <= conv1_bias_array[0];\
					added_1[94] <= conv1_bias_array[0];\
					added_1[95] <= conv1_bias_array[0];\
					added_1[96] <= conv1_bias_array[0];\
					added_1[97] <= conv1_bias_array[0];\
					added_1[98] <= conv1_bias_array[0];\
					added_1[99] <= conv1_bias_array[0];\
					added_1[100] <= conv1_bias_array[0];\
					added_1[101] <= conv1_bias_array[0];\
					added_1[102] <= conv1_bias_array[0];\
					added_1[103] <= conv1_bias_array[0];\
					added_1[104] <= conv1_bias_array[0];\
					added_1[105] <= conv1_bias_array[0];\
					added_1[106] <= conv1_bias_array[0];\
					added_1[107] <= conv1_bias_array[0];\
					added_1[108] <= conv1_bias_array[0];\
					added_1[109] <= conv1_bias_array[0];\
					added_1[110] <= conv1_bias_array[0];\
					added_1[111] <= conv1_bias_array[0];\
                end\
                else if(cnt2<8'd6) begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_1[110] <= product_result[110];\
					added_1[111] <= product_result[111];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
					added_2[110] <= add_result[110];\
					added_2[111] <= add_result[111];\
                end\
                else begin\
                    added_2[0] <= 18'd0;\
                    added_2[1] <= 18'd0;\
                    added_2[2] <= 18'd0;\
                    added_2[3] <= 18'd0;\
                    added_2[4] <= 18'd0;\
                    added_2[5] <= 18'd0;\
                    added_2[6] <= 18'd0;\
                    added_2[7] <= 18'd0;\
                    added_2[8] <= 18'd0;\
                    added_2[9] <= 18'd0;\
                    added_2[10] <= 18'd0;\
                    added_2[11] <= 18'd0;\
                    added_2[12] <= 18'd0;\
                    added_2[13] <= 18'd0;\
                    added_2[14] <= 18'd0;\
                    added_2[15] <= 18'd0;\
                    added_2[16] <= 18'd0;\
                    added_2[17] <= 18'd0;\
                    added_2[18] <= 18'd0;\
                    added_2[19] <= 18'd0;\
                    added_2[20] <= 18'd0;\
                    added_2[21] <= 18'd0;\
                    added_2[22] <= 18'd0;\
                    added_2[23] <= 18'd0;\
                    added_2[24] <= 18'd0;\
                    added_2[25] <= 18'd0;\
                    added_2[26] <= 18'd0;\
                    added_2[27] <= 18'd0;\
                    added_2[28] <= 18'd0;\
                    added_2[29] <= 18'd0;\
                    added_2[30] <= 18'd0;\
                    added_2[31] <= 18'd0;\
                    added_2[32] <= 18'd0;\
                    added_2[33] <= 18'd0;\
                    added_2[34] <= 18'd0;\
                    added_2[35] <= 18'd0;\
                    added_2[36] <= 18'd0;\
                    added_2[37] <= 18'd0;\
                    added_2[38] <= 18'd0;\
                    added_2[39] <= 18'd0;\
                    added_2[40] <= 18'd0;\
                    added_2[41] <= 18'd0;\
                    added_2[42] <= 18'd0;\
                    added_2[43] <= 18'd0;\
                    added_2[44] <= 18'd0;\
                    added_2[45] <= 18'd0;\
                    added_2[46] <= 18'd0;\
                    added_2[47] <= 18'd0;\
                    added_2[48] <= 18'd0;\
                    added_2[49] <= 18'd0;\
                    added_2[50] <= 18'd0;\
                    added_2[51] <= 18'd0;\
                    added_2[52] <= 18'd0;\
                    added_2[53] <= 18'd0;\
                    added_2[54] <= 18'd0;\
                    added_2[55] <= 18'd0;\
                    added_2[56] <= 18'd0;\
                    added_2[57] <= 18'd0;\
                    added_2[58] <= 18'd0;\
                    added_2[59] <= 18'd0;\
                    added_2[60] <= 18'd0;\
                    added_2[61] <= 18'd0;\
                    added_2[62] <= 18'd0;\
                    added_2[63] <= 18'd0;\
                    added_2[64] <= 18'd0;\
                    added_2[65] <= 18'd0;\
                    added_2[66] <= 18'd0;\
                    added_2[67] <= 18'd0;\
                    added_2[68] <= 18'd0;\
                    added_2[69] <= 18'd0;\
                    added_2[70] <= 18'd0;\
                    added_2[71] <= 18'd0;\
                    added_2[72] <= 18'd0;\
                    added_2[73] <= 18'd0;\
                    added_2[74] <= 18'd0;\
                    added_2[75] <= 18'd0;\
                    added_2[76] <= 18'd0;\
                    added_2[77] <= 18'd0;\
                    added_2[78] <= 18'd0;\
                    added_2[79] <= 18'd0;\
                    added_2[80] <= 18'd0;\
                    added_2[81] <= 18'd0;\
                    added_2[82] <= 18'd0;\
                    added_2[83] <= 18'd0;\
                    added_2[84] <= 18'd0;\
                    added_2[85] <= 18'd0;\
                    added_2[86] <= 18'd0;\
                    added_2[87] <= 18'd0;\
                    added_2[88] <= 18'd0;\
                    added_2[89] <= 18'd0;\
                    added_2[90] <= 18'd0;\
                    added_2[91] <= 18'd0;\
                    added_2[92] <= 18'd0;\
                    added_2[93] <= 18'd0;\
                    added_2[94] <= 18'd0;\
                    added_2[95] <= 18'd0;\
                    added_2[96] <= 18'd0;\
                    added_2[97] <= 18'd0;\
                    added_2[98] <= 18'd0;\
                    added_2[99] <= 18'd0;\
                    added_2[100] <= 18'd0;\
                    added_2[101] <= 18'd0;\
                    added_2[102] <= 18'd0;\
                    added_2[103] <= 18'd0;\
                    added_2[104] <= 18'd0;\
                    added_2[105] <= 18'd0;\
                    added_2[106] <= 18'd0;\
                    added_2[107] <= 18'd0;\
                    added_2[108] <= 18'd0;\
                    added_2[109] <= 18'd0;\
                    added_2[110] <= 18'd0;\
                    added_2[111] <= 18'd0;\
                end\
            end\
            CONV1_2_1,CONV1_2_2,CONV1_2_3,CONV1_2_4,CONV1_2_5,CONV1_2_6,CONV1_2_7:begin \
                if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[0] <= conv1_bias_array[1];\
					added_1[1] <= conv1_bias_array[1];\
					added_1[2] <= conv1_bias_array[1];\
					added_1[3] <= conv1_bias_array[1];\
					added_1[4] <= conv1_bias_array[1];\
					added_1[5] <= conv1_bias_array[1];\
					added_1[6] <= conv1_bias_array[1];\
					added_1[7] <= conv1_bias_array[1];\
					added_1[8] <= conv1_bias_array[1];\
					added_1[9] <= conv1_bias_array[1];\
					added_1[10] <= conv1_bias_array[1];\
					added_1[11] <= conv1_bias_array[1];\
					added_1[12] <= conv1_bias_array[1];\
					added_1[13] <= conv1_bias_array[1];\
					added_1[14] <= conv1_bias_array[1];\
					added_1[15] <= conv1_bias_array[1];\
					added_1[16] <= conv1_bias_array[1];\
					added_1[17] <= conv1_bias_array[1];\
					added_1[18] <= conv1_bias_array[1];\
					added_1[19] <= conv1_bias_array[1];\
					added_1[20] <= conv1_bias_array[1];\
					added_1[21] <= conv1_bias_array[1];\
					added_1[22] <= conv1_bias_array[1];\
					added_1[23] <= conv1_bias_array[1];\
					added_1[24] <= conv1_bias_array[1];\
					added_1[25] <= conv1_bias_array[1];\
					added_1[26] <= conv1_bias_array[1];\
					added_1[27] <= conv1_bias_array[1];\
					added_1[28] <= conv1_bias_array[1];\
					added_1[29] <= conv1_bias_array[1];\
					added_1[30] <= conv1_bias_array[1];\
					added_1[31] <= conv1_bias_array[1];\
					added_1[32] <= conv1_bias_array[1];\
					added_1[33] <= conv1_bias_array[1];\
					added_1[34] <= conv1_bias_array[1];\
					added_1[35] <= conv1_bias_array[1];\
					added_1[36] <= conv1_bias_array[1];\
					added_1[37] <= conv1_bias_array[1];\
					added_1[38] <= conv1_bias_array[1];\
					added_1[39] <= conv1_bias_array[1];\
					added_1[40] <= conv1_bias_array[1];\
					added_1[41] <= conv1_bias_array[1];\
					added_1[42] <= conv1_bias_array[1];\
					added_1[43] <= conv1_bias_array[1];\
					added_1[44] <= conv1_bias_array[1];\
					added_1[45] <= conv1_bias_array[1];\
					added_1[46] <= conv1_bias_array[1];\
					added_1[47] <= conv1_bias_array[1];\
					added_1[48] <= conv1_bias_array[1];\
					added_1[49] <= conv1_bias_array[1];\
					added_1[50] <= conv1_bias_array[1];\
					added_1[51] <= conv1_bias_array[1];\
					added_1[52] <= conv1_bias_array[1];\
					added_1[53] <= conv1_bias_array[1];\
					added_1[54] <= conv1_bias_array[1];\
					added_1[55] <= conv1_bias_array[1];\
					added_1[56] <= conv1_bias_array[1];\
					added_1[57] <= conv1_bias_array[1];\
					added_1[58] <= conv1_bias_array[1];\
					added_1[59] <= conv1_bias_array[1];\
					added_1[60] <= conv1_bias_array[1];\
					added_1[61] <= conv1_bias_array[1];\
					added_1[62] <= conv1_bias_array[1];\
					added_1[63] <= conv1_bias_array[1];\
					added_1[64] <= conv1_bias_array[1];\
					added_1[65] <= conv1_bias_array[1];\
					added_1[66] <= conv1_bias_array[1];\
					added_1[67] <= conv1_bias_array[1];\
					added_1[68] <= conv1_bias_array[1];\
					added_1[69] <= conv1_bias_array[1];\
					added_1[70] <= conv1_bias_array[1];\
					added_1[71] <= conv1_bias_array[1];\
					added_1[72] <= conv1_bias_array[1];\
					added_1[73] <= conv1_bias_array[1];\
					added_1[74] <= conv1_bias_array[1];\
					added_1[75] <= conv1_bias_array[1];\
					added_1[76] <= conv1_bias_array[1];\
					added_1[77] <= conv1_bias_array[1];\
					added_1[78] <= conv1_bias_array[1];\
					added_1[79] <= conv1_bias_array[1];\
					added_1[80] <= conv1_bias_array[1];\
					added_1[81] <= conv1_bias_array[1];\
					added_1[82] <= conv1_bias_array[1];\
					added_1[83] <= conv1_bias_array[1];\
					added_1[84] <= conv1_bias_array[1];\
					added_1[85] <= conv1_bias_array[1];\
					added_1[86] <= conv1_bias_array[1];\
					added_1[87] <= conv1_bias_array[1];\
					added_1[88] <= conv1_bias_array[1];\
					added_1[89] <= conv1_bias_array[1];\
					added_1[90] <= conv1_bias_array[1];\
					added_1[91] <= conv1_bias_array[1];\
					added_1[92] <= conv1_bias_array[1];\
					added_1[93] <= conv1_bias_array[1];\
					added_1[94] <= conv1_bias_array[1];\
					added_1[95] <= conv1_bias_array[1];\
					added_1[96] <= conv1_bias_array[1];\
					added_1[97] <= conv1_bias_array[1];\
					added_1[98] <= conv1_bias_array[1];\
					added_1[99] <= conv1_bias_array[1];\
					added_1[100] <= conv1_bias_array[1];\
					added_1[101] <= conv1_bias_array[1];\
					added_1[102] <= conv1_bias_array[1];\
					added_1[103] <= conv1_bias_array[1];\
					added_1[104] <= conv1_bias_array[1];\
					added_1[105] <= conv1_bias_array[1];\
					added_1[106] <= conv1_bias_array[1];\
					added_1[107] <= conv1_bias_array[1];\
					added_1[108] <= conv1_bias_array[1];\
					added_1[109] <= conv1_bias_array[1];\
					added_1[110] <= conv1_bias_array[1];\
					added_1[111] <= conv1_bias_array[1];\
                end\
                else if(cnt2<8'd6) begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_1[110] <= product_result[110];\
					added_1[111] <= product_result[111];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
					added_2[110] <= add_result[110];\
					added_2[111] <= add_result[111];\
                end\
                else begin\
                    added_2[0] <= 18'd0;\
                    added_2[1] <= 18'd0;\
                    added_2[2] <= 18'd0;\
                    added_2[3] <= 18'd0;\
                    added_2[4] <= 18'd0;\
                    added_2[5] <= 18'd0;\
                    added_2[6] <= 18'd0;\
                    added_2[7] <= 18'd0;\
                    added_2[8] <= 18'd0;\
                    added_2[9] <= 18'd0;\
                    added_2[10] <= 18'd0;\
                    added_2[11] <= 18'd0;\
                    added_2[12] <= 18'd0;\
                    added_2[13] <= 18'd0;\
                    added_2[14] <= 18'd0;\
                    added_2[15] <= 18'd0;\
                    added_2[16] <= 18'd0;\
                    added_2[17] <= 18'd0;\
                    added_2[18] <= 18'd0;\
                    added_2[19] <= 18'd0;\
                    added_2[20] <= 18'd0;\
                    added_2[21] <= 18'd0;\
                    added_2[22] <= 18'd0;\
                    added_2[23] <= 18'd0;\
                    added_2[24] <= 18'd0;\
                    added_2[25] <= 18'd0;\
                    added_2[26] <= 18'd0;\
                    added_2[27] <= 18'd0;\
                    added_2[28] <= 18'd0;\
                    added_2[29] <= 18'd0;\
                    added_2[30] <= 18'd0;\
                    added_2[31] <= 18'd0;\
                    added_2[32] <= 18'd0;\
                    added_2[33] <= 18'd0;\
                    added_2[34] <= 18'd0;\
                    added_2[35] <= 18'd0;\
                    added_2[36] <= 18'd0;\
                    added_2[37] <= 18'd0;\
                    added_2[38] <= 18'd0;\
                    added_2[39] <= 18'd0;\
                    added_2[40] <= 18'd0;\
                    added_2[41] <= 18'd0;\
                    added_2[42] <= 18'd0;\
                    added_2[43] <= 18'd0;\
                    added_2[44] <= 18'd0;\
                    added_2[45] <= 18'd0;\
                    added_2[46] <= 18'd0;\
                    added_2[47] <= 18'd0;\
                    added_2[48] <= 18'd0;\
                    added_2[49] <= 18'd0;\
                    added_2[50] <= 18'd0;\
                    added_2[51] <= 18'd0;\
                    added_2[52] <= 18'd0;\
                    added_2[53] <= 18'd0;\
                    added_2[54] <= 18'd0;\
                    added_2[55] <= 18'd0;\
                    added_2[56] <= 18'd0;\
                    added_2[57] <= 18'd0;\
                    added_2[58] <= 18'd0;\
                    added_2[59] <= 18'd0;\
                    added_2[60] <= 18'd0;\
                    added_2[61] <= 18'd0;\
                    added_2[62] <= 18'd0;\
                    added_2[63] <= 18'd0;\
                    added_2[64] <= 18'd0;\
                    added_2[65] <= 18'd0;\
                    added_2[66] <= 18'd0;\
                    added_2[67] <= 18'd0;\
                    added_2[68] <= 18'd0;\
                    added_2[69] <= 18'd0;\
                    added_2[70] <= 18'd0;\
                    added_2[71] <= 18'd0;\
                    added_2[72] <= 18'd0;\
                    added_2[73] <= 18'd0;\
                    added_2[74] <= 18'd0;\
                    added_2[75] <= 18'd0;\
                    added_2[76] <= 18'd0;\
                    added_2[77] <= 18'd0;\
                    added_2[78] <= 18'd0;\
                    added_2[79] <= 18'd0;\
                    added_2[80] <= 18'd0;\
                    added_2[81] <= 18'd0;\
                    added_2[82] <= 18'd0;\
                    added_2[83] <= 18'd0;\
                    added_2[84] <= 18'd0;\
                    added_2[85] <= 18'd0;\
                    added_2[86] <= 18'd0;\
                    added_2[87] <= 18'd0;\
                    added_2[88] <= 18'd0;\
                    added_2[89] <= 18'd0;\
                    added_2[90] <= 18'd0;\
                    added_2[91] <= 18'd0;\
                    added_2[92] <= 18'd0;\
                    added_2[93] <= 18'd0;\
                    added_2[94] <= 18'd0;\
                    added_2[95] <= 18'd0;\
                    added_2[96] <= 18'd0;\
                    added_2[97] <= 18'd0;\
                    added_2[98] <= 18'd0;\
                    added_2[99] <= 18'd0;\
                    added_2[100] <= 18'd0;\
                    added_2[101] <= 18'd0;\
                    added_2[102] <= 18'd0;\
                    added_2[103] <= 18'd0;\
                    added_2[104] <= 18'd0;\
                    added_2[105] <= 18'd0;\
                    added_2[106] <= 18'd0;\
                    added_2[107] <= 18'd0;\
                    added_2[108] <= 18'd0;\
                    added_2[109] <= 18'd0;\
                    added_2[110] <= 18'd0;\
                    added_2[111] <= 18'd0;\
                end\
            end\
            CONV1_3_1,CONV1_3_2,CONV1_3_3,CONV1_3_4,CONV1_3_5,CONV1_3_6,CONV1_3_7:begin \
                if((cnt1==8'd0)&(cnt2==8'd0))begin\
					added_1[0] <= conv1_bias_array[2];\
					added_1[1] <= conv1_bias_array[2];\
					added_1[2] <= conv1_bias_array[2];\
					added_1[3] <= conv1_bias_array[2];\
					added_1[4] <= conv1_bias_array[2];\
					added_1[5] <= conv1_bias_array[2];\
					added_1[6] <= conv1_bias_array[2];\
					added_1[7] <= conv1_bias_array[2];\
					added_1[8] <= conv1_bias_array[2];\
					added_1[9] <= conv1_bias_array[2];\
					added_1[10] <= conv1_bias_array[2];\
					added_1[11] <= conv1_bias_array[2];\
					added_1[12] <= conv1_bias_array[2];\
					added_1[13] <= conv1_bias_array[2];\
					added_1[14] <= conv1_bias_array[2];\
					added_1[15] <= conv1_bias_array[2];\
					added_1[16] <= conv1_bias_array[2];\
					added_1[17] <= conv1_bias_array[2];\
					added_1[18] <= conv1_bias_array[2];\
					added_1[19] <= conv1_bias_array[2];\
					added_1[20] <= conv1_bias_array[2];\
					added_1[21] <= conv1_bias_array[2];\
					added_1[22] <= conv1_bias_array[2];\
					added_1[23] <= conv1_bias_array[2];\
					added_1[24] <= conv1_bias_array[2];\
					added_1[25] <= conv1_bias_array[2];\
					added_1[26] <= conv1_bias_array[2];\
					added_1[27] <= conv1_bias_array[2];\
					added_1[28] <= conv1_bias_array[2];\
					added_1[29] <= conv1_bias_array[2];\
					added_1[30] <= conv1_bias_array[2];\
					added_1[31] <= conv1_bias_array[2];\
					added_1[32] <= conv1_bias_array[2];\
					added_1[33] <= conv1_bias_array[2];\
					added_1[34] <= conv1_bias_array[2];\
					added_1[35] <= conv1_bias_array[2];\
					added_1[36] <= conv1_bias_array[2];\
					added_1[37] <= conv1_bias_array[2];\
					added_1[38] <= conv1_bias_array[2];\
					added_1[39] <= conv1_bias_array[2];\
					added_1[40] <= conv1_bias_array[2];\
					added_1[41] <= conv1_bias_array[2];\
					added_1[42] <= conv1_bias_array[2];\
					added_1[43] <= conv1_bias_array[2];\
					added_1[44] <= conv1_bias_array[2];\
					added_1[45] <= conv1_bias_array[2];\
					added_1[46] <= conv1_bias_array[2];\
					added_1[47] <= conv1_bias_array[2];\
					added_1[48] <= conv1_bias_array[2];\
					added_1[49] <= conv1_bias_array[2];\
					added_1[50] <= conv1_bias_array[2];\
					added_1[51] <= conv1_bias_array[2];\
					added_1[52] <= conv1_bias_array[2];\
					added_1[53] <= conv1_bias_array[2];\
					added_1[54] <= conv1_bias_array[2];\
					added_1[55] <= conv1_bias_array[2];\
					added_1[56] <= conv1_bias_array[2];\
					added_1[57] <= conv1_bias_array[2];\
					added_1[58] <= conv1_bias_array[2];\
					added_1[59] <= conv1_bias_array[2];\
					added_1[60] <= conv1_bias_array[2];\
					added_1[61] <= conv1_bias_array[2];\
					added_1[62] <= conv1_bias_array[2];\
					added_1[63] <= conv1_bias_array[2];\
					added_1[64] <= conv1_bias_array[2];\
					added_1[65] <= conv1_bias_array[2];\
					added_1[66] <= conv1_bias_array[2];\
					added_1[67] <= conv1_bias_array[2];\
					added_1[68] <= conv1_bias_array[2];\
					added_1[69] <= conv1_bias_array[2];\
					added_1[70] <= conv1_bias_array[2];\
					added_1[71] <= conv1_bias_array[2];\
					added_1[72] <= conv1_bias_array[2];\
					added_1[73] <= conv1_bias_array[2];\
					added_1[74] <= conv1_bias_array[2];\
					added_1[75] <= conv1_bias_array[2];\
					added_1[76] <= conv1_bias_array[2];\
					added_1[77] <= conv1_bias_array[2];\
					added_1[78] <= conv1_bias_array[2];\
					added_1[79] <= conv1_bias_array[2];\
					added_1[80] <= conv1_bias_array[2];\
					added_1[81] <= conv1_bias_array[2];\
					added_1[82] <= conv1_bias_array[2];\
					added_1[83] <= conv1_bias_array[2];\
					added_1[84] <= conv1_bias_array[2];\
					added_1[85] <= conv1_bias_array[2];\
					added_1[86] <= conv1_bias_array[2];\
					added_1[87] <= conv1_bias_array[2];\
					added_1[88] <= conv1_bias_array[2];\
					added_1[89] <= conv1_bias_array[2];\
					added_1[90] <= conv1_bias_array[2];\
					added_1[91] <= conv1_bias_array[2];\
					added_1[92] <= conv1_bias_array[2];\
					added_1[93] <= conv1_bias_array[2];\
					added_1[94] <= conv1_bias_array[2];\
					added_1[95] <= conv1_bias_array[2];\
					added_1[96] <= conv1_bias_array[2];\
					added_1[97] <= conv1_bias_array[2];\
					added_1[98] <= conv1_bias_array[2];\
					added_1[99] <= conv1_bias_array[2];\
					added_1[100] <= conv1_bias_array[2];\
					added_1[101] <= conv1_bias_array[2];\
					added_1[102] <= conv1_bias_array[2];\
					added_1[103] <= conv1_bias_array[2];\
					added_1[104] <= conv1_bias_array[2];\
					added_1[105] <= conv1_bias_array[2];\
					added_1[106] <= conv1_bias_array[2];\
					added_1[107] <= conv1_bias_array[2];\
					added_1[108] <= conv1_bias_array[2];\
					added_1[109] <= conv1_bias_array[2];\
					added_1[110] <= conv1_bias_array[2];\
					added_1[111] <= conv1_bias_array[2];\
                end\
                else if(cnt2<8'd6) begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_1[110] <= product_result[110];\
					added_1[111] <= product_result[111];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
					added_2[110] <= add_result[110];\
					added_2[111] <= add_result[111];\
                end\
                else begin\
                    added_2[0] <= 18'd0;\
                    added_2[1] <= 18'd0;\
                    added_2[2] <= 18'd0;\
                    added_2[3] <= 18'd0;\
                    added_2[4] <= 18'd0;\
                    added_2[5] <= 18'd0;\
                    added_2[6] <= 18'd0;\
                    added_2[7] <= 18'd0;\
                    added_2[8] <= 18'd0;\
                    added_2[9] <= 18'd0;\
                    added_2[10] <= 18'd0;\
                    added_2[11] <= 18'd0;\
                    added_2[12] <= 18'd0;\
                    added_2[13] <= 18'd0;\
                    added_2[14] <= 18'd0;\
                    added_2[15] <= 18'd0;\
                    added_2[16] <= 18'd0;\
                    added_2[17] <= 18'd0;\
                    added_2[18] <= 18'd0;\
                    added_2[19] <= 18'd0;\
                    added_2[20] <= 18'd0;\
                    added_2[21] <= 18'd0;\
                    added_2[22] <= 18'd0;\
                    added_2[23] <= 18'd0;\
                    added_2[24] <= 18'd0;\
                    added_2[25] <= 18'd0;\
                    added_2[26] <= 18'd0;\
                    added_2[27] <= 18'd0;\
                    added_2[28] <= 18'd0;\
                    added_2[29] <= 18'd0;\
                    added_2[30] <= 18'd0;\
                    added_2[31] <= 18'd0;\
                    added_2[32] <= 18'd0;\
                    added_2[33] <= 18'd0;\
                    added_2[34] <= 18'd0;\
                    added_2[35] <= 18'd0;\
                    added_2[36] <= 18'd0;\
                    added_2[37] <= 18'd0;\
                    added_2[38] <= 18'd0;\
                    added_2[39] <= 18'd0;\
                    added_2[40] <= 18'd0;\
                    added_2[41] <= 18'd0;\
                    added_2[42] <= 18'd0;\
                    added_2[43] <= 18'd0;\
                    added_2[44] <= 18'd0;\
                    added_2[45] <= 18'd0;\
                    added_2[46] <= 18'd0;\
                    added_2[47] <= 18'd0;\
                    added_2[48] <= 18'd0;\
                    added_2[49] <= 18'd0;\
                    added_2[50] <= 18'd0;\
                    added_2[51] <= 18'd0;\
                    added_2[52] <= 18'd0;\
                    added_2[53] <= 18'd0;\
                    added_2[54] <= 18'd0;\
                    added_2[55] <= 18'd0;\
                    added_2[56] <= 18'd0;\
                    added_2[57] <= 18'd0;\
                    added_2[58] <= 18'd0;\
                    added_2[59] <= 18'd0;\
                    added_2[60] <= 18'd0;\
                    added_2[61] <= 18'd0;\
                    added_2[62] <= 18'd0;\
                    added_2[63] <= 18'd0;\
                    added_2[64] <= 18'd0;\
                    added_2[65] <= 18'd0;\
                    added_2[66] <= 18'd0;\
                    added_2[67] <= 18'd0;\
                    added_2[68] <= 18'd0;\
                    added_2[69] <= 18'd0;\
                    added_2[70] <= 18'd0;\
                    added_2[71] <= 18'd0;\
                    added_2[72] <= 18'd0;\
                    added_2[73] <= 18'd0;\
                    added_2[74] <= 18'd0;\
                    added_2[75] <= 18'd0;\
                    added_2[76] <= 18'd0;\
                    added_2[77] <= 18'd0;\
                    added_2[78] <= 18'd0;\
                    added_2[79] <= 18'd0;\
                    added_2[80] <= 18'd0;\
                    added_2[81] <= 18'd0;\
                    added_2[82] <= 18'd0;\
                    added_2[83] <= 18'd0;\
                    added_2[84] <= 18'd0;\
                    added_2[85] <= 18'd0;\
                    added_2[86] <= 18'd0;\
                    added_2[87] <= 18'd0;\
                    added_2[88] <= 18'd0;\
                    added_2[89] <= 18'd0;\
                    added_2[90] <= 18'd0;\
                    added_2[91] <= 18'd0;\
                    added_2[92] <= 18'd0;\
                    added_2[93] <= 18'd0;\
                    added_2[94] <= 18'd0;\
                    added_2[95] <= 18'd0;\
                    added_2[96] <= 18'd0;\
                    added_2[97] <= 18'd0;\
                    added_2[98] <= 18'd0;\
                    added_2[99] <= 18'd0;\
                    added_2[100] <= 18'd0;\
                    added_2[101] <= 18'd0;\
                    added_2[102] <= 18'd0;\
                    added_2[103] <= 18'd0;\
                    added_2[104] <= 18'd0;\
                    added_2[105] <= 18'd0;\
                    added_2[106] <= 18'd0;\
                    added_2[107] <= 18'd0;\
                    added_2[108] <= 18'd0;\
                    added_2[109] <= 18'd0;\
                    added_2[110] <= 18'd0;\
                    added_2[111] <= 18'd0;\
                end\
            end\
            CONV1_4_1,CONV1_4_2,CONV1_4_3,CONV1_4_4,CONV1_4_5,CONV1_4_6,CONV1_4_7:begin \
                if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[0] <= conv1_bias_array[3];\
					added_1[1] <= conv1_bias_array[3];\
					added_1[2] <= conv1_bias_array[3];\
					added_1[3] <= conv1_bias_array[3];\
					added_1[4] <= conv1_bias_array[3];\
					added_1[5] <= conv1_bias_array[3];\
					added_1[6] <= conv1_bias_array[3];\
					added_1[7] <= conv1_bias_array[3];\
					added_1[8] <= conv1_bias_array[3];\
					added_1[9] <= conv1_bias_array[3];\
					added_1[10] <= conv1_bias_array[3];\
					added_1[11] <= conv1_bias_array[3];\
					added_1[12] <= conv1_bias_array[3];\
					added_1[13] <= conv1_bias_array[3];\
					added_1[14] <= conv1_bias_array[3];\
					added_1[15] <= conv1_bias_array[3];\
					added_1[16] <= conv1_bias_array[3];\
					added_1[17] <= conv1_bias_array[3];\
					added_1[18] <= conv1_bias_array[3];\
					added_1[19] <= conv1_bias_array[3];\
					added_1[20] <= conv1_bias_array[3];\
					added_1[21] <= conv1_bias_array[3];\
					added_1[22] <= conv1_bias_array[3];\
					added_1[23] <= conv1_bias_array[3];\
					added_1[24] <= conv1_bias_array[3];\
					added_1[25] <= conv1_bias_array[3];\
					added_1[26] <= conv1_bias_array[3];\
					added_1[27] <= conv1_bias_array[3];\
					added_1[28] <= conv1_bias_array[3];\
					added_1[29] <= conv1_bias_array[3];\
					added_1[30] <= conv1_bias_array[3];\
					added_1[31] <= conv1_bias_array[3];\
					added_1[32] <= conv1_bias_array[3];\
					added_1[33] <= conv1_bias_array[3];\
					added_1[34] <= conv1_bias_array[3];\
					added_1[35] <= conv1_bias_array[3];\
					added_1[36] <= conv1_bias_array[3];\
					added_1[37] <= conv1_bias_array[3];\
					added_1[38] <= conv1_bias_array[3];\
					added_1[39] <= conv1_bias_array[3];\
					added_1[40] <= conv1_bias_array[3];\
					added_1[41] <= conv1_bias_array[3];\
					added_1[42] <= conv1_bias_array[3];\
					added_1[43] <= conv1_bias_array[3];\
					added_1[44] <= conv1_bias_array[3];\
					added_1[45] <= conv1_bias_array[3];\
					added_1[46] <= conv1_bias_array[3];\
					added_1[47] <= conv1_bias_array[3];\
					added_1[48] <= conv1_bias_array[3];\
					added_1[49] <= conv1_bias_array[3];\
					added_1[50] <= conv1_bias_array[3];\
					added_1[51] <= conv1_bias_array[3];\
					added_1[52] <= conv1_bias_array[3];\
					added_1[53] <= conv1_bias_array[3];\
					added_1[54] <= conv1_bias_array[3];\
					added_1[55] <= conv1_bias_array[3];\
					added_1[56] <= conv1_bias_array[3];\
					added_1[57] <= conv1_bias_array[3];\
					added_1[58] <= conv1_bias_array[3];\
					added_1[59] <= conv1_bias_array[3];\
					added_1[60] <= conv1_bias_array[3];\
					added_1[61] <= conv1_bias_array[3];\
					added_1[62] <= conv1_bias_array[3];\
					added_1[63] <= conv1_bias_array[3];\
					added_1[64] <= conv1_bias_array[3];\
					added_1[65] <= conv1_bias_array[3];\
					added_1[66] <= conv1_bias_array[3];\
					added_1[67] <= conv1_bias_array[3];\
					added_1[68] <= conv1_bias_array[3];\
					added_1[69] <= conv1_bias_array[3];\
					added_1[70] <= conv1_bias_array[3];\
					added_1[71] <= conv1_bias_array[3];\
					added_1[72] <= conv1_bias_array[3];\
					added_1[73] <= conv1_bias_array[3];\
					added_1[74] <= conv1_bias_array[3];\
					added_1[75] <= conv1_bias_array[3];\
					added_1[76] <= conv1_bias_array[3];\
					added_1[77] <= conv1_bias_array[3];\
					added_1[78] <= conv1_bias_array[3];\
					added_1[79] <= conv1_bias_array[3];\
					added_1[80] <= conv1_bias_array[3];\
					added_1[81] <= conv1_bias_array[3];\
					added_1[82] <= conv1_bias_array[3];\
					added_1[83] <= conv1_bias_array[3];\
					added_1[84] <= conv1_bias_array[3];\
					added_1[85] <= conv1_bias_array[3];\
					added_1[86] <= conv1_bias_array[3];\
					added_1[87] <= conv1_bias_array[3];\
					added_1[88] <= conv1_bias_array[3];\
					added_1[89] <= conv1_bias_array[3];\
					added_1[90] <= conv1_bias_array[3];\
					added_1[91] <= conv1_bias_array[3];\
					added_1[92] <= conv1_bias_array[3];\
					added_1[93] <= conv1_bias_array[3];\
					added_1[94] <= conv1_bias_array[3];\
					added_1[95] <= conv1_bias_array[3];\
					added_1[96] <= conv1_bias_array[3];\
					added_1[97] <= conv1_bias_array[3];\
					added_1[98] <= conv1_bias_array[3];\
					added_1[99] <= conv1_bias_array[3];\
					added_1[100] <= conv1_bias_array[3];\
					added_1[101] <= conv1_bias_array[3];\
					added_1[102] <= conv1_bias_array[3];\
					added_1[103] <= conv1_bias_array[3];\
					added_1[104] <= conv1_bias_array[3];\
					added_1[105] <= conv1_bias_array[3];\
					added_1[106] <= conv1_bias_array[3];\
					added_1[107] <= conv1_bias_array[3];\
					added_1[108] <= conv1_bias_array[3];\
					added_1[109] <= conv1_bias_array[3];\
					added_1[110] <= conv1_bias_array[3];\
					added_1[111] <= conv1_bias_array[3];\
                end\
                else if(cnt2<8'd6) begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_1[110] <= product_result[110];\
					added_1[111] <= product_result[111];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
					added_2[110] <= add_result[110];\
					added_2[111] <= add_result[111];\
                end\
                else begin\
                    added_2[0] <= 18'd0;\
                    added_2[1] <= 18'd0;\
                    added_2[2] <= 18'd0;\
                    added_2[3] <= 18'd0;\
                    added_2[4] <= 18'd0;\
                    added_2[5] <= 18'd0;\
                    added_2[6] <= 18'd0;\
                    added_2[7] <= 18'd0;\
                    added_2[8] <= 18'd0;\
                    added_2[9] <= 18'd0;\
                    added_2[10] <= 18'd0;\
                    added_2[11] <= 18'd0;\
                    added_2[12] <= 18'd0;\
                    added_2[13] <= 18'd0;\
                    added_2[14] <= 18'd0;\
                    added_2[15] <= 18'd0;\
                    added_2[16] <= 18'd0;\
                    added_2[17] <= 18'd0;\
                    added_2[18] <= 18'd0;\
                    added_2[19] <= 18'd0;\
                    added_2[20] <= 18'd0;\
                    added_2[21] <= 18'd0;\
                    added_2[22] <= 18'd0;\
                    added_2[23] <= 18'd0;\
                    added_2[24] <= 18'd0;\
                    added_2[25] <= 18'd0;\
                    added_2[26] <= 18'd0;\
                    added_2[27] <= 18'd0;\
                    added_2[28] <= 18'd0;\
                    added_2[29] <= 18'd0;\
                    added_2[30] <= 18'd0;\
                    added_2[31] <= 18'd0;\
                    added_2[32] <= 18'd0;\
                    added_2[33] <= 18'd0;\
                    added_2[34] <= 18'd0;\
                    added_2[35] <= 18'd0;\
                    added_2[36] <= 18'd0;\
                    added_2[37] <= 18'd0;\
                    added_2[38] <= 18'd0;\
                    added_2[39] <= 18'd0;\
                    added_2[40] <= 18'd0;\
                    added_2[41] <= 18'd0;\
                    added_2[42] <= 18'd0;\
                    added_2[43] <= 18'd0;\
                    added_2[44] <= 18'd0;\
                    added_2[45] <= 18'd0;\
                    added_2[46] <= 18'd0;\
                    added_2[47] <= 18'd0;\
                    added_2[48] <= 18'd0;\
                    added_2[49] <= 18'd0;\
                    added_2[50] <= 18'd0;\
                    added_2[51] <= 18'd0;\
                    added_2[52] <= 18'd0;\
                    added_2[53] <= 18'd0;\
                    added_2[54] <= 18'd0;\
                    added_2[55] <= 18'd0;\
                    added_2[56] <= 18'd0;\
                    added_2[57] <= 18'd0;\
                    added_2[58] <= 18'd0;\
                    added_2[59] <= 18'd0;\
                    added_2[60] <= 18'd0;\
                    added_2[61] <= 18'd0;\
                    added_2[62] <= 18'd0;\
                    added_2[63] <= 18'd0;\
                    added_2[64] <= 18'd0;\
                    added_2[65] <= 18'd0;\
                    added_2[66] <= 18'd0;\
                    added_2[67] <= 18'd0;\
                    added_2[68] <= 18'd0;\
                    added_2[69] <= 18'd0;\
                    added_2[70] <= 18'd0;\
                    added_2[71] <= 18'd0;\
                    added_2[72] <= 18'd0;\
                    added_2[73] <= 18'd0;\
                    added_2[74] <= 18'd0;\
                    added_2[75] <= 18'd0;\
                    added_2[76] <= 18'd0;\
                    added_2[77] <= 18'd0;\
                    added_2[78] <= 18'd0;\
                    added_2[79] <= 18'd0;\
                    added_2[80] <= 18'd0;\
                    added_2[81] <= 18'd0;\
                    added_2[82] <= 18'd0;\
                    added_2[83] <= 18'd0;\
                    added_2[84] <= 18'd0;\
                    added_2[85] <= 18'd0;\
                    added_2[86] <= 18'd0;\
                    added_2[87] <= 18'd0;\
                    added_2[88] <= 18'd0;\
                    added_2[89] <= 18'd0;\
                    added_2[90] <= 18'd0;\
                    added_2[91] <= 18'd0;\
                    added_2[92] <= 18'd0;\
                    added_2[93] <= 18'd0;\
                    added_2[94] <= 18'd0;\
                    added_2[95] <= 18'd0;\
                    added_2[96] <= 18'd0;\
                    added_2[97] <= 18'd0;\
                    added_2[98] <= 18'd0;\
                    added_2[99] <= 18'd0;\
                    added_2[100] <= 18'd0;\
                    added_2[101] <= 18'd0;\
                    added_2[102] <= 18'd0;\
                    added_2[103] <= 18'd0;\
                    added_2[104] <= 18'd0;\
                    added_2[105] <= 18'd0;\
                    added_2[106] <= 18'd0;\
                    added_2[107] <= 18'd0;\
                    added_2[108] <= 18'd0;\
                    added_2[109] <= 18'd0;\
                    added_2[110] <= 18'd0;\
                    added_2[111] <= 18'd0;\
                end\
            end\
            CONV1_5_1,CONV1_5_2,CONV1_5_3,CONV1_5_4,CONV1_5_5,CONV1_5_6,CONV1_5_7:begin \
                if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[0] <= conv1_bias_array[4];\
					added_1[1] <= conv1_bias_array[4];\
					added_1[2] <= conv1_bias_array[4];\
					added_1[3] <= conv1_bias_array[4];\
					added_1[4] <= conv1_bias_array[4];\
					added_1[5] <= conv1_bias_array[4];\
					added_1[6] <= conv1_bias_array[4];\
					added_1[7] <= conv1_bias_array[4];\
					added_1[8] <= conv1_bias_array[4];\
					added_1[9] <= conv1_bias_array[4];\
					added_1[10] <= conv1_bias_array[4];\
					added_1[11] <= conv1_bias_array[4];\
					added_1[12] <= conv1_bias_array[4];\
					added_1[13] <= conv1_bias_array[4];\
					added_1[14] <= conv1_bias_array[4];\
					added_1[15] <= conv1_bias_array[4];\
					added_1[16] <= conv1_bias_array[4];\
					added_1[17] <= conv1_bias_array[4];\
					added_1[18] <= conv1_bias_array[4];\
					added_1[19] <= conv1_bias_array[4];\
					added_1[20] <= conv1_bias_array[4];\
					added_1[21] <= conv1_bias_array[4];\
					added_1[22] <= conv1_bias_array[4];\
					added_1[23] <= conv1_bias_array[4];\
					added_1[24] <= conv1_bias_array[4];\
					added_1[25] <= conv1_bias_array[4];\
					added_1[26] <= conv1_bias_array[4];\
					added_1[27] <= conv1_bias_array[4];\
					added_1[28] <= conv1_bias_array[4];\
					added_1[29] <= conv1_bias_array[4];\
					added_1[30] <= conv1_bias_array[4];\
					added_1[31] <= conv1_bias_array[4];\
					added_1[32] <= conv1_bias_array[4];\
					added_1[33] <= conv1_bias_array[4];\
					added_1[34] <= conv1_bias_array[4];\
					added_1[35] <= conv1_bias_array[4];\
					added_1[36] <= conv1_bias_array[4];\
					added_1[37] <= conv1_bias_array[4];\
					added_1[38] <= conv1_bias_array[4];\
					added_1[39] <= conv1_bias_array[4];\
					added_1[40] <= conv1_bias_array[4];\
					added_1[41] <= conv1_bias_array[4];\
					added_1[42] <= conv1_bias_array[4];\
					added_1[43] <= conv1_bias_array[4];\
					added_1[44] <= conv1_bias_array[4];\
					added_1[45] <= conv1_bias_array[4];\
					added_1[46] <= conv1_bias_array[4];\
					added_1[47] <= conv1_bias_array[4];\
					added_1[48] <= conv1_bias_array[4];\
					added_1[49] <= conv1_bias_array[4];\
					added_1[50] <= conv1_bias_array[4];\
					added_1[51] <= conv1_bias_array[4];\
					added_1[52] <= conv1_bias_array[4];\
					added_1[53] <= conv1_bias_array[4];\
					added_1[54] <= conv1_bias_array[4];\
					added_1[55] <= conv1_bias_array[4];\
					added_1[56] <= conv1_bias_array[4];\
					added_1[57] <= conv1_bias_array[4];\
					added_1[58] <= conv1_bias_array[4];\
					added_1[59] <= conv1_bias_array[4];\
					added_1[60] <= conv1_bias_array[4];\
					added_1[61] <= conv1_bias_array[4];\
					added_1[62] <= conv1_bias_array[4];\
					added_1[63] <= conv1_bias_array[4];\
					added_1[64] <= conv1_bias_array[4];\
					added_1[65] <= conv1_bias_array[4];\
					added_1[66] <= conv1_bias_array[4];\
					added_1[67] <= conv1_bias_array[4];\
					added_1[68] <= conv1_bias_array[4];\
					added_1[69] <= conv1_bias_array[4];\
					added_1[70] <= conv1_bias_array[4];\
					added_1[71] <= conv1_bias_array[4];\
					added_1[72] <= conv1_bias_array[4];\
					added_1[73] <= conv1_bias_array[4];\
					added_1[74] <= conv1_bias_array[4];\
					added_1[75] <= conv1_bias_array[4];\
					added_1[76] <= conv1_bias_array[4];\
					added_1[77] <= conv1_bias_array[4];\
					added_1[78] <= conv1_bias_array[4];\
					added_1[79] <= conv1_bias_array[4];\
					added_1[80] <= conv1_bias_array[4];\
					added_1[81] <= conv1_bias_array[4];\
					added_1[82] <= conv1_bias_array[4];\
					added_1[83] <= conv1_bias_array[4];\
					added_1[84] <= conv1_bias_array[4];\
					added_1[85] <= conv1_bias_array[4];\
					added_1[86] <= conv1_bias_array[4];\
					added_1[87] <= conv1_bias_array[4];\
					added_1[88] <= conv1_bias_array[4];\
					added_1[89] <= conv1_bias_array[4];\
					added_1[90] <= conv1_bias_array[4];\
					added_1[91] <= conv1_bias_array[4];\
					added_1[92] <= conv1_bias_array[4];\
					added_1[93] <= conv1_bias_array[4];\
					added_1[94] <= conv1_bias_array[4];\
					added_1[95] <= conv1_bias_array[4];\
					added_1[96] <= conv1_bias_array[4];\
					added_1[97] <= conv1_bias_array[4];\
					added_1[98] <= conv1_bias_array[4];\
					added_1[99] <= conv1_bias_array[4];\
					added_1[100] <= conv1_bias_array[4];\
					added_1[101] <= conv1_bias_array[4];\
					added_1[102] <= conv1_bias_array[4];\
					added_1[103] <= conv1_bias_array[4];\
					added_1[104] <= conv1_bias_array[4];\
					added_1[105] <= conv1_bias_array[4];\
					added_1[106] <= conv1_bias_array[4];\
					added_1[107] <= conv1_bias_array[4];\
					added_1[108] <= conv1_bias_array[4];\
					added_1[109] <= conv1_bias_array[4];\
					added_1[110] <= conv1_bias_array[4];\
					added_1[111] <= conv1_bias_array[4];\
                end\
                else if(cnt2<8'd6) begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_1[110] <= product_result[110];\
					added_1[111] <= product_result[111];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
					added_2[110] <= add_result[110];\
					added_2[111] <= add_result[111];\
                end\
                else begin\
                    added_2[0] <= 18'd0;\
                    added_2[1] <= 18'd0;\
                    added_2[2] <= 18'd0;\
                    added_2[3] <= 18'd0;\
                    added_2[4] <= 18'd0;\
                    added_2[5] <= 18'd0;\
                    added_2[6] <= 18'd0;\
                    added_2[7] <= 18'd0;\
                    added_2[8] <= 18'd0;\
                    added_2[9] <= 18'd0;\
                    added_2[10] <= 18'd0;\
                    added_2[11] <= 18'd0;\
                    added_2[12] <= 18'd0;\
                    added_2[13] <= 18'd0;\
                    added_2[14] <= 18'd0;\
                    added_2[15] <= 18'd0;\
                    added_2[16] <= 18'd0;\
                    added_2[17] <= 18'd0;\
                    added_2[18] <= 18'd0;\
                    added_2[19] <= 18'd0;\
                    added_2[20] <= 18'd0;\
                    added_2[21] <= 18'd0;\
                    added_2[22] <= 18'd0;\
                    added_2[23] <= 18'd0;\
                    added_2[24] <= 18'd0;\
                    added_2[25] <= 18'd0;\
                    added_2[26] <= 18'd0;\
                    added_2[27] <= 18'd0;\
                    added_2[28] <= 18'd0;\
                    added_2[29] <= 18'd0;\
                    added_2[30] <= 18'd0;\
                    added_2[31] <= 18'd0;\
                    added_2[32] <= 18'd0;\
                    added_2[33] <= 18'd0;\
                    added_2[34] <= 18'd0;\
                    added_2[35] <= 18'd0;\
                    added_2[36] <= 18'd0;\
                    added_2[37] <= 18'd0;\
                    added_2[38] <= 18'd0;\
                    added_2[39] <= 18'd0;\
                    added_2[40] <= 18'd0;\
                    added_2[41] <= 18'd0;\
                    added_2[42] <= 18'd0;\
                    added_2[43] <= 18'd0;\
                    added_2[44] <= 18'd0;\
                    added_2[45] <= 18'd0;\
                    added_2[46] <= 18'd0;\
                    added_2[47] <= 18'd0;\
                    added_2[48] <= 18'd0;\
                    added_2[49] <= 18'd0;\
                    added_2[50] <= 18'd0;\
                    added_2[51] <= 18'd0;\
                    added_2[52] <= 18'd0;\
                    added_2[53] <= 18'd0;\
                    added_2[54] <= 18'd0;\
                    added_2[55] <= 18'd0;\
                    added_2[56] <= 18'd0;\
                    added_2[57] <= 18'd0;\
                    added_2[58] <= 18'd0;\
                    added_2[59] <= 18'd0;\
                    added_2[60] <= 18'd0;\
                    added_2[61] <= 18'd0;\
                    added_2[62] <= 18'd0;\
                    added_2[63] <= 18'd0;\
                    added_2[64] <= 18'd0;\
                    added_2[65] <= 18'd0;\
                    added_2[66] <= 18'd0;\
                    added_2[67] <= 18'd0;\
                    added_2[68] <= 18'd0;\
                    added_2[69] <= 18'd0;\
                    added_2[70] <= 18'd0;\
                    added_2[71] <= 18'd0;\
                    added_2[72] <= 18'd0;\
                    added_2[73] <= 18'd0;\
                    added_2[74] <= 18'd0;\
                    added_2[75] <= 18'd0;\
                    added_2[76] <= 18'd0;\
                    added_2[77] <= 18'd0;\
                    added_2[78] <= 18'd0;\
                    added_2[79] <= 18'd0;\
                    added_2[80] <= 18'd0;\
                    added_2[81] <= 18'd0;\
                    added_2[82] <= 18'd0;\
                    added_2[83] <= 18'd0;\
                    added_2[84] <= 18'd0;\
                    added_2[85] <= 18'd0;\
                    added_2[86] <= 18'd0;\
                    added_2[87] <= 18'd0;\
                    added_2[88] <= 18'd0;\
                    added_2[89] <= 18'd0;\
                    added_2[90] <= 18'd0;\
                    added_2[91] <= 18'd0;\
                    added_2[92] <= 18'd0;\
                    added_2[93] <= 18'd0;\
                    added_2[94] <= 18'd0;\
                    added_2[95] <= 18'd0;\
                    added_2[96] <= 18'd0;\
                    added_2[97] <= 18'd0;\
                    added_2[98] <= 18'd0;\
                    added_2[99] <= 18'd0;\
                    added_2[100] <= 18'd0;\
                    added_2[101] <= 18'd0;\
                    added_2[102] <= 18'd0;\
                    added_2[103] <= 18'd0;\
                    added_2[104] <= 18'd0;\
                    added_2[105] <= 18'd0;\
                    added_2[106] <= 18'd0;\
                    added_2[107] <= 18'd0;\
                    added_2[108] <= 18'd0;\
                    added_2[109] <= 18'd0;\
                    added_2[110] <= 18'd0;\
                    added_2[111] <= 18'd0;\
                end\
            end\
            CONV1_6_1,CONV1_6_2,CONV1_6_3,CONV1_6_4,CONV1_6_5,CONV1_6_6,CONV1_6_7:begin \
                if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[0] <= conv1_bias_array[5];\
					added_1[1] <= conv1_bias_array[5];\
					added_1[2] <= conv1_bias_array[5];\
					added_1[3] <= conv1_bias_array[5];\
					added_1[4] <= conv1_bias_array[5];\
					added_1[5] <= conv1_bias_array[5];\
					added_1[6] <= conv1_bias_array[5];\
					added_1[7] <= conv1_bias_array[5];\
					added_1[8] <= conv1_bias_array[5];\
					added_1[9] <= conv1_bias_array[5];\
					added_1[10] <= conv1_bias_array[5];\
					added_1[11] <= conv1_bias_array[5];\
					added_1[12] <= conv1_bias_array[5];\
					added_1[13] <= conv1_bias_array[5];\
					added_1[14] <= conv1_bias_array[5];\
					added_1[15] <= conv1_bias_array[5];\
					added_1[16] <= conv1_bias_array[5];\
					added_1[17] <= conv1_bias_array[5];\
					added_1[18] <= conv1_bias_array[5];\
					added_1[19] <= conv1_bias_array[5];\
					added_1[20] <= conv1_bias_array[5];\
					added_1[21] <= conv1_bias_array[5];\
					added_1[22] <= conv1_bias_array[5];\
					added_1[23] <= conv1_bias_array[5];\
					added_1[24] <= conv1_bias_array[5];\
					added_1[25] <= conv1_bias_array[5];\
					added_1[26] <= conv1_bias_array[5];\
					added_1[27] <= conv1_bias_array[5];\
					added_1[28] <= conv1_bias_array[5];\
					added_1[29] <= conv1_bias_array[5];\
					added_1[30] <= conv1_bias_array[5];\
					added_1[31] <= conv1_bias_array[5];\
					added_1[32] <= conv1_bias_array[5];\
					added_1[33] <= conv1_bias_array[5];\
					added_1[34] <= conv1_bias_array[5];\
					added_1[35] <= conv1_bias_array[5];\
					added_1[36] <= conv1_bias_array[5];\
					added_1[37] <= conv1_bias_array[5];\
					added_1[38] <= conv1_bias_array[5];\
					added_1[39] <= conv1_bias_array[5];\
					added_1[40] <= conv1_bias_array[5];\
					added_1[41] <= conv1_bias_array[5];\
					added_1[42] <= conv1_bias_array[5];\
					added_1[43] <= conv1_bias_array[5];\
					added_1[44] <= conv1_bias_array[5];\
					added_1[45] <= conv1_bias_array[5];\
					added_1[46] <= conv1_bias_array[5];\
					added_1[47] <= conv1_bias_array[5];\
					added_1[48] <= conv1_bias_array[5];\
					added_1[49] <= conv1_bias_array[5];\
					added_1[50] <= conv1_bias_array[5];\
					added_1[51] <= conv1_bias_array[5];\
					added_1[52] <= conv1_bias_array[5];\
					added_1[53] <= conv1_bias_array[5];\
					added_1[54] <= conv1_bias_array[5];\
					added_1[55] <= conv1_bias_array[5];\
					added_1[56] <= conv1_bias_array[5];\
					added_1[57] <= conv1_bias_array[5];\
					added_1[58] <= conv1_bias_array[5];\
					added_1[59] <= conv1_bias_array[5];\
					added_1[60] <= conv1_bias_array[5];\
					added_1[61] <= conv1_bias_array[5];\
					added_1[62] <= conv1_bias_array[5];\
					added_1[63] <= conv1_bias_array[5];\
					added_1[64] <= conv1_bias_array[5];\
					added_1[65] <= conv1_bias_array[5];\
					added_1[66] <= conv1_bias_array[5];\
					added_1[67] <= conv1_bias_array[5];\
					added_1[68] <= conv1_bias_array[5];\
					added_1[69] <= conv1_bias_array[5];\
					added_1[70] <= conv1_bias_array[5];\
					added_1[71] <= conv1_bias_array[5];\
					added_1[72] <= conv1_bias_array[5];\
					added_1[73] <= conv1_bias_array[5];\
					added_1[74] <= conv1_bias_array[5];\
					added_1[75] <= conv1_bias_array[5];\
					added_1[76] <= conv1_bias_array[5];\
					added_1[77] <= conv1_bias_array[5];\
					added_1[78] <= conv1_bias_array[5];\
					added_1[79] <= conv1_bias_array[5];\
					added_1[80] <= conv1_bias_array[5];\
					added_1[81] <= conv1_bias_array[5];\
					added_1[82] <= conv1_bias_array[5];\
					added_1[83] <= conv1_bias_array[5];\
					added_1[84] <= conv1_bias_array[5];\
					added_1[85] <= conv1_bias_array[5];\
					added_1[86] <= conv1_bias_array[5];\
					added_1[87] <= conv1_bias_array[5];\
					added_1[88] <= conv1_bias_array[5];\
					added_1[89] <= conv1_bias_array[5];\
					added_1[90] <= conv1_bias_array[5];\
					added_1[91] <= conv1_bias_array[5];\
					added_1[92] <= conv1_bias_array[5];\
					added_1[93] <= conv1_bias_array[5];\
					added_1[94] <= conv1_bias_array[5];\
					added_1[95] <= conv1_bias_array[5];\
					added_1[96] <= conv1_bias_array[5];\
					added_1[97] <= conv1_bias_array[5];\
					added_1[98] <= conv1_bias_array[5];\
					added_1[99] <= conv1_bias_array[5];\
					added_1[100] <= conv1_bias_array[5];\
					added_1[101] <= conv1_bias_array[5];\
					added_1[102] <= conv1_bias_array[5];\
					added_1[103] <= conv1_bias_array[5];\
					added_1[104] <= conv1_bias_array[5];\
					added_1[105] <= conv1_bias_array[5];\
					added_1[106] <= conv1_bias_array[5];\
					added_1[107] <= conv1_bias_array[5];\
					added_1[108] <= conv1_bias_array[5];\
					added_1[109] <= conv1_bias_array[5];\
					added_1[110] <= conv1_bias_array[5];\
					added_1[111] <= conv1_bias_array[5];\
                end\
                else if(cnt2<8'd6) begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_1[110] <= product_result[110];\
					added_1[111] <= product_result[111];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
					added_2[110] <= add_result[110];\
					added_2[111] <= add_result[111];\
                end\
                else begin\
                    added_2[0] <= 18'd0;\
                    added_2[1] <= 18'd0;\
                    added_2[2] <= 18'd0;\
                    added_2[3] <= 18'd0;\
                    added_2[4] <= 18'd0;\
                    added_2[5] <= 18'd0;\
                    added_2[6] <= 18'd0;\
                    added_2[7] <= 18'd0;\
                    added_2[8] <= 18'd0;\
                    added_2[9] <= 18'd0;\
                    added_2[10] <= 18'd0;\
                    added_2[11] <= 18'd0;\
                    added_2[12] <= 18'd0;\
                    added_2[13] <= 18'd0;\
                    added_2[14] <= 18'd0;\
                    added_2[15] <= 18'd0;\
                    added_2[16] <= 18'd0;\
                    added_2[17] <= 18'd0;\
                    added_2[18] <= 18'd0;\
                    added_2[19] <= 18'd0;\
                    added_2[20] <= 18'd0;\
                    added_2[21] <= 18'd0;\
                    added_2[22] <= 18'd0;\
                    added_2[23] <= 18'd0;\
                    added_2[24] <= 18'd0;\
                    added_2[25] <= 18'd0;\
                    added_2[26] <= 18'd0;\
                    added_2[27] <= 18'd0;\
                    added_2[28] <= 18'd0;\
                    added_2[29] <= 18'd0;\
                    added_2[30] <= 18'd0;\
                    added_2[31] <= 18'd0;\
                    added_2[32] <= 18'd0;\
                    added_2[33] <= 18'd0;\
                    added_2[34] <= 18'd0;\
                    added_2[35] <= 18'd0;\
                    added_2[36] <= 18'd0;\
                    added_2[37] <= 18'd0;\
                    added_2[38] <= 18'd0;\
                    added_2[39] <= 18'd0;\
                    added_2[40] <= 18'd0;\
                    added_2[41] <= 18'd0;\
                    added_2[42] <= 18'd0;\
                    added_2[43] <= 18'd0;\
                    added_2[44] <= 18'd0;\
                    added_2[45] <= 18'd0;\
                    added_2[46] <= 18'd0;\
                    added_2[47] <= 18'd0;\
                    added_2[48] <= 18'd0;\
                    added_2[49] <= 18'd0;\
                    added_2[50] <= 18'd0;\
                    added_2[51] <= 18'd0;\
                    added_2[52] <= 18'd0;\
                    added_2[53] <= 18'd0;\
                    added_2[54] <= 18'd0;\
                    added_2[55] <= 18'd0;\
                    added_2[56] <= 18'd0;\
                    added_2[57] <= 18'd0;\
                    added_2[58] <= 18'd0;\
                    added_2[59] <= 18'd0;\
                    added_2[60] <= 18'd0;\
                    added_2[61] <= 18'd0;\
                    added_2[62] <= 18'd0;\
                    added_2[63] <= 18'd0;\
                    added_2[64] <= 18'd0;\
                    added_2[65] <= 18'd0;\
                    added_2[66] <= 18'd0;\
                    added_2[67] <= 18'd0;\
                    added_2[68] <= 18'd0;\
                    added_2[69] <= 18'd0;\
                    added_2[70] <= 18'd0;\
                    added_2[71] <= 18'd0;\
                    added_2[72] <= 18'd0;\
                    added_2[73] <= 18'd0;\
                    added_2[74] <= 18'd0;\
                    added_2[75] <= 18'd0;\
                    added_2[76] <= 18'd0;\
                    added_2[77] <= 18'd0;\
                    added_2[78] <= 18'd0;\
                    added_2[79] <= 18'd0;\
                    added_2[80] <= 18'd0;\
                    added_2[81] <= 18'd0;\
                    added_2[82] <= 18'd0;\
                    added_2[83] <= 18'd0;\
                    added_2[84] <= 18'd0;\
                    added_2[85] <= 18'd0;\
                    added_2[86] <= 18'd0;\
                    added_2[87] <= 18'd0;\
                    added_2[88] <= 18'd0;\
                    added_2[89] <= 18'd0;\
                    added_2[90] <= 18'd0;\
                    added_2[91] <= 18'd0;\
                    added_2[92] <= 18'd0;\
                    added_2[93] <= 18'd0;\
                    added_2[94] <= 18'd0;\
                    added_2[95] <= 18'd0;\
                    added_2[96] <= 18'd0;\
                    added_2[97] <= 18'd0;\
                    added_2[98] <= 18'd0;\
                    added_2[99] <= 18'd0;\
                    added_2[100] <= 18'd0;\
                    added_2[101] <= 18'd0;\
                    added_2[102] <= 18'd0;\
                    added_2[103] <= 18'd0;\
                    added_2[104] <= 18'd0;\
                    added_2[105] <= 18'd0;\
                    added_2[106] <= 18'd0;\
                    added_2[107] <= 18'd0;\
                    added_2[108] <= 18'd0;\
                    added_2[109] <= 18'd0;\
                    added_2[110] <= 18'd0;\
                    added_2[111] <= 18'd0;\
                end\
            end\
            CONV2_1_1:begin\
				if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[ 0] <= conv2_bias_array[0];\
					added_1[ 1] <= conv2_bias_array[0];\
					added_1[ 2] <= conv2_bias_array[0];\
					added_1[ 3] <= conv2_bias_array[0];\
					added_1[ 4] <= conv2_bias_array[0];\
					added_1[ 5] <= conv2_bias_array[0];\
					added_1[ 6] <= conv2_bias_array[0];\
					added_1[ 7] <= conv2_bias_array[0];\
					added_1[ 8] <= conv2_bias_array[0];\
					added_1[ 9] <= conv2_bias_array[0];\
					added_1[10] <= conv2_bias_array[0];\
					added_1[11] <= conv2_bias_array[0];\
					added_1[12] <= conv2_bias_array[0];\
					added_1[13] <= conv2_bias_array[0];\
					added_1[14] <= conv2_bias_array[0];\
					added_1[15] <= conv2_bias_array[0];\
					added_1[16] <= conv2_bias_array[0];\
					added_1[17] <= conv2_bias_array[0];\
					added_1[18] <= conv2_bias_array[0];\
					added_1[19] <= conv2_bias_array[0];\
					added_1[20] <= conv2_bias_array[0];\
					added_1[21] <= conv2_bias_array[0];\
					added_1[22] <= conv2_bias_array[0];\
					added_1[23] <= conv2_bias_array[0];\
					added_1[24] <= conv2_bias_array[0];\
					added_1[25] <= conv2_bias_array[0];\
					added_1[26] <= conv2_bias_array[0];\
					added_1[27] <= conv2_bias_array[0];\
					added_1[28] <= conv2_bias_array[0];\
					added_1[29] <= conv2_bias_array[0];\
					added_1[30] <= conv2_bias_array[0];\
					added_1[31] <= conv2_bias_array[0];\
					added_1[32] <= conv2_bias_array[0];\
					added_1[33] <= conv2_bias_array[0];\
					added_1[34] <= conv2_bias_array[0];\
					added_1[35] <= conv2_bias_array[0];\
					added_1[36] <= conv2_bias_array[0];\
					added_1[37] <= conv2_bias_array[0];\
					added_1[38] <= conv2_bias_array[0];\
					added_1[39] <= conv2_bias_array[0];\
					added_1[40] <= conv2_bias_array[0];\
					added_1[41] <= conv2_bias_array[0];\
					added_1[42] <= conv2_bias_array[0];\
					added_1[43] <= conv2_bias_array[0];\
					added_1[44] <= conv2_bias_array[0];\
					added_1[45] <= conv2_bias_array[0];\
					added_1[46] <= conv2_bias_array[0];\
					added_1[47] <= conv2_bias_array[0];\
					added_1[48] <= conv2_bias_array[0];\
					added_1[49] <= conv2_bias_array[0];\
					added_1[50] <= conv2_bias_array[0];\
					added_1[51] <= conv2_bias_array[0];\
					added_1[52] <= conv2_bias_array[0];\
					added_1[53] <= conv2_bias_array[0];\
					added_1[54] <= conv2_bias_array[0];\
					added_1[55] <= conv2_bias_array[0];\
					added_1[56] <= conv2_bias_array[0];\
					added_1[57] <= conv2_bias_array[0];\
					added_1[58] <= conv2_bias_array[0];\
					added_1[59] <= conv2_bias_array[0];\
					added_1[60] <= conv2_bias_array[0];\
					added_1[61] <= conv2_bias_array[0];\
					added_1[62] <= conv2_bias_array[0];\
					added_1[63] <= conv2_bias_array[0];\
					added_1[64] <= conv2_bias_array[0];\
					added_1[65] <= conv2_bias_array[0];\
					added_1[66] <= conv2_bias_array[0];\
					added_1[67] <= conv2_bias_array[0];\
					added_1[68] <= conv2_bias_array[0];\
					added_1[69] <= conv2_bias_array[0];\
					added_1[70] <= conv2_bias_array[0];\
					added_1[71] <= conv2_bias_array[0];\
					added_1[72] <= conv2_bias_array[0];\
					added_1[73] <= conv2_bias_array[0];\
					added_1[74] <= conv2_bias_array[0];\
					added_1[75] <= conv2_bias_array[0];\
					added_1[76] <= conv2_bias_array[0];\
					added_1[77] <= conv2_bias_array[0];\
					added_1[78] <= conv2_bias_array[0];\
					added_1[79] <= conv2_bias_array[0];\
					added_1[80] <= conv2_bias_array[0];\
					added_1[81] <= conv2_bias_array[0];\
					added_1[82] <= conv2_bias_array[0];\
					added_1[83] <= conv2_bias_array[0];\
					added_1[84] <= conv2_bias_array[0];\
					added_1[85] <= conv2_bias_array[0];\
					added_1[86] <= conv2_bias_array[0];\
					added_1[87] <= conv2_bias_array[0];\
					added_1[88] <= conv2_bias_array[0];\
					added_1[89] <= conv2_bias_array[0];\
					added_1[90] <= conv2_bias_array[0];\
					added_1[91] <= conv2_bias_array[0];\
					added_1[92] <= conv2_bias_array[0];\
					added_1[93] <= conv2_bias_array[0];\
					added_1[94] <= conv2_bias_array[0];\
					added_1[95] <= conv2_bias_array[0];\
					added_1[96] <= conv2_bias_array[0];\
					added_1[97] <= conv2_bias_array[0];\
					added_1[98] <= conv2_bias_array[0];\
					added_1[99] <= conv2_bias_array[0];\
				end\
				else begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
				end\
			end\
			CONV2_2_1:begin\
				if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[ 0] <= conv2_bias_array[1];\
					added_1[ 1] <= conv2_bias_array[1];\
					added_1[ 2] <= conv2_bias_array[1];\
					added_1[ 3] <= conv2_bias_array[1];\
					added_1[ 4] <= conv2_bias_array[1];\
					added_1[ 5] <= conv2_bias_array[1];\
					added_1[ 6] <= conv2_bias_array[1];\
					added_1[ 7] <= conv2_bias_array[1];\
					added_1[ 8] <= conv2_bias_array[1];\
					added_1[ 9] <= conv2_bias_array[1];\
					added_1[10] <= conv2_bias_array[1];\
					added_1[11] <= conv2_bias_array[1];\
					added_1[12] <= conv2_bias_array[1];\
					added_1[13] <= conv2_bias_array[1];\
					added_1[14] <= conv2_bias_array[1];\
					added_1[15] <= conv2_bias_array[1];\
					added_1[16] <= conv2_bias_array[1];\
					added_1[17] <= conv2_bias_array[1];\
					added_1[18] <= conv2_bias_array[1];\
					added_1[19] <= conv2_bias_array[1];\
					added_1[20] <= conv2_bias_array[1];\
					added_1[21] <= conv2_bias_array[1];\
					added_1[22] <= conv2_bias_array[1];\
					added_1[23] <= conv2_bias_array[1];\
					added_1[24] <= conv2_bias_array[1];\
					added_1[25] <= conv2_bias_array[1];\
					added_1[26] <= conv2_bias_array[1];\
					added_1[27] <= conv2_bias_array[1];\
					added_1[28] <= conv2_bias_array[1];\
					added_1[29] <= conv2_bias_array[1];\
					added_1[30] <= conv2_bias_array[1];\
					added_1[31] <= conv2_bias_array[1];\
					added_1[32] <= conv2_bias_array[1];\
					added_1[33] <= conv2_bias_array[1];\
					added_1[34] <= conv2_bias_array[1];\
					added_1[35] <= conv2_bias_array[1];\
					added_1[36] <= conv2_bias_array[1];\
					added_1[37] <= conv2_bias_array[1];\
					added_1[38] <= conv2_bias_array[1];\
					added_1[39] <= conv2_bias_array[1];\
					added_1[40] <= conv2_bias_array[1];\
					added_1[41] <= conv2_bias_array[1];\
					added_1[42] <= conv2_bias_array[1];\
					added_1[43] <= conv2_bias_array[1];\
					added_1[44] <= conv2_bias_array[1];\
					added_1[45] <= conv2_bias_array[1];\
					added_1[46] <= conv2_bias_array[1];\
					added_1[47] <= conv2_bias_array[1];\
					added_1[48] <= conv2_bias_array[1];\
					added_1[49] <= conv2_bias_array[1];\
					added_1[50] <= conv2_bias_array[1];\
					added_1[51] <= conv2_bias_array[1];\
					added_1[52] <= conv2_bias_array[1];\
					added_1[53] <= conv2_bias_array[1];\
					added_1[54] <= conv2_bias_array[1];\
					added_1[55] <= conv2_bias_array[1];\
					added_1[56] <= conv2_bias_array[1];\
					added_1[57] <= conv2_bias_array[1];\
					added_1[58] <= conv2_bias_array[1];\
					added_1[59] <= conv2_bias_array[1];\
					added_1[60] <= conv2_bias_array[1];\
					added_1[61] <= conv2_bias_array[1];\
					added_1[62] <= conv2_bias_array[1];\
					added_1[63] <= conv2_bias_array[1];\
					added_1[64] <= conv2_bias_array[1];\
					added_1[65] <= conv2_bias_array[1];\
					added_1[66] <= conv2_bias_array[1];\
					added_1[67] <= conv2_bias_array[1];\
					added_1[68] <= conv2_bias_array[1];\
					added_1[69] <= conv2_bias_array[1];\
					added_1[70] <= conv2_bias_array[1];\
					added_1[71] <= conv2_bias_array[1];\
					added_1[72] <= conv2_bias_array[1];\
					added_1[73] <= conv2_bias_array[1];\
					added_1[74] <= conv2_bias_array[1];\
					added_1[75] <= conv2_bias_array[1];\
					added_1[76] <= conv2_bias_array[1];\
					added_1[77] <= conv2_bias_array[1];\
					added_1[78] <= conv2_bias_array[1];\
					added_1[79] <= conv2_bias_array[1];\
					added_1[80] <= conv2_bias_array[1];\
					added_1[81] <= conv2_bias_array[1];\
					added_1[82] <= conv2_bias_array[1];\
					added_1[83] <= conv2_bias_array[1];\
					added_1[84] <= conv2_bias_array[1];\
					added_1[85] <= conv2_bias_array[1];\
					added_1[86] <= conv2_bias_array[1];\
					added_1[87] <= conv2_bias_array[1];\
					added_1[88] <= conv2_bias_array[1];\
					added_1[89] <= conv2_bias_array[1];\
					added_1[90] <= conv2_bias_array[1];\
					added_1[91] <= conv2_bias_array[1];\
					added_1[92] <= conv2_bias_array[1];\
					added_1[93] <= conv2_bias_array[1];\
					added_1[94] <= conv2_bias_array[1];\
					added_1[95] <= conv2_bias_array[1];\
					added_1[96] <= conv2_bias_array[1];\
					added_1[97] <= conv2_bias_array[1];\
					added_1[98] <= conv2_bias_array[1];\
					added_1[99] <= conv2_bias_array[1];\
				end\
				else begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
				end\
			end\
            CONV2_3_1:begin\
				if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[ 0] <= conv2_bias_array[2];\
					added_1[ 1] <= conv2_bias_array[2];\
					added_1[ 2] <= conv2_bias_array[2];\
					added_1[ 3] <= conv2_bias_array[2];\
					added_1[ 4] <= conv2_bias_array[2];\
					added_1[ 5] <= conv2_bias_array[2];\
					added_1[ 6] <= conv2_bias_array[2];\
					added_1[ 7] <= conv2_bias_array[2];\
					added_1[ 8] <= conv2_bias_array[2];\
					added_1[ 9] <= conv2_bias_array[2];\
					added_1[10] <= conv2_bias_array[2];\
					added_1[11] <= conv2_bias_array[2];\
					added_1[12] <= conv2_bias_array[2];\
					added_1[13] <= conv2_bias_array[2];\
					added_1[14] <= conv2_bias_array[2];\
					added_1[15] <= conv2_bias_array[2];\
					added_1[16] <= conv2_bias_array[2];\
					added_1[17] <= conv2_bias_array[2];\
					added_1[18] <= conv2_bias_array[2];\
					added_1[19] <= conv2_bias_array[2];\
					added_1[20] <= conv2_bias_array[2];\
					added_1[21] <= conv2_bias_array[2];\
					added_1[22] <= conv2_bias_array[2];\
					added_1[23] <= conv2_bias_array[2];\
					added_1[24] <= conv2_bias_array[2];\
					added_1[25] <= conv2_bias_array[2];\
					added_1[26] <= conv2_bias_array[2];\
					added_1[27] <= conv2_bias_array[2];\
					added_1[28] <= conv2_bias_array[2];\
					added_1[29] <= conv2_bias_array[2];\
					added_1[30] <= conv2_bias_array[2];\
					added_1[31] <= conv2_bias_array[2];\
					added_1[32] <= conv2_bias_array[2];\
					added_1[33] <= conv2_bias_array[2];\
					added_1[34] <= conv2_bias_array[2];\
					added_1[35] <= conv2_bias_array[2];\
					added_1[36] <= conv2_bias_array[2];\
					added_1[37] <= conv2_bias_array[2];\
					added_1[38] <= conv2_bias_array[2];\
					added_1[39] <= conv2_bias_array[2];\
					added_1[40] <= conv2_bias_array[2];\
					added_1[41] <= conv2_bias_array[2];\
					added_1[42] <= conv2_bias_array[2];\
					added_1[43] <= conv2_bias_array[2];\
					added_1[44] <= conv2_bias_array[2];\
					added_1[45] <= conv2_bias_array[2];\
					added_1[46] <= conv2_bias_array[2];\
					added_1[47] <= conv2_bias_array[2];\
					added_1[48] <= conv2_bias_array[2];\
					added_1[49] <= conv2_bias_array[2];\
					added_1[50] <= conv2_bias_array[2];\
					added_1[51] <= conv2_bias_array[2];\
					added_1[52] <= conv2_bias_array[2];\
					added_1[53] <= conv2_bias_array[2];\
					added_1[54] <= conv2_bias_array[2];\
					added_1[55] <= conv2_bias_array[2];\
					added_1[56] <= conv2_bias_array[2];\
					added_1[57] <= conv2_bias_array[2];\
					added_1[58] <= conv2_bias_array[2];\
					added_1[59] <= conv2_bias_array[2];\
					added_1[60] <= conv2_bias_array[2];\
					added_1[61] <= conv2_bias_array[2];\
					added_1[62] <= conv2_bias_array[2];\
					added_1[63] <= conv2_bias_array[2];\
					added_1[64] <= conv2_bias_array[2];\
					added_1[65] <= conv2_bias_array[2];\
					added_1[66] <= conv2_bias_array[2];\
					added_1[67] <= conv2_bias_array[2];\
					added_1[68] <= conv2_bias_array[2];\
					added_1[69] <= conv2_bias_array[2];\
					added_1[70] <= conv2_bias_array[2];\
					added_1[71] <= conv2_bias_array[2];\
					added_1[72] <= conv2_bias_array[2];\
					added_1[73] <= conv2_bias_array[2];\
					added_1[74] <= conv2_bias_array[2];\
					added_1[75] <= conv2_bias_array[2];\
					added_1[76] <= conv2_bias_array[2];\
					added_1[77] <= conv2_bias_array[2];\
					added_1[78] <= conv2_bias_array[2];\
					added_1[79] <= conv2_bias_array[2];\
					added_1[80] <= conv2_bias_array[2];\
					added_1[81] <= conv2_bias_array[2];\
					added_1[82] <= conv2_bias_array[2];\
					added_1[83] <= conv2_bias_array[2];\
					added_1[84] <= conv2_bias_array[2];\
					added_1[85] <= conv2_bias_array[2];\
					added_1[86] <= conv2_bias_array[2];\
					added_1[87] <= conv2_bias_array[2];\
					added_1[88] <= conv2_bias_array[2];\
					added_1[89] <= conv2_bias_array[2];\
					added_1[90] <= conv2_bias_array[2];\
					added_1[91] <= conv2_bias_array[2];\
					added_1[92] <= conv2_bias_array[2];\
					added_1[93] <= conv2_bias_array[2];\
					added_1[94] <= conv2_bias_array[2];\
					added_1[95] <= conv2_bias_array[2];\
					added_1[96] <= conv2_bias_array[2];\
					added_1[97] <= conv2_bias_array[2];\
					added_1[98] <= conv2_bias_array[2];\
					added_1[99] <= conv2_bias_array[2];\
				end\
				else begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
				end\
			end\
            CONV2_4_1:begin\
				if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[ 0] <= conv2_bias_array[3];\
					added_1[ 1] <= conv2_bias_array[3];\
					added_1[ 2] <= conv2_bias_array[3];\
					added_1[ 3] <= conv2_bias_array[3];\
					added_1[ 4] <= conv2_bias_array[3];\
					added_1[ 5] <= conv2_bias_array[3];\
					added_1[ 6] <= conv2_bias_array[3];\
					added_1[ 7] <= conv2_bias_array[3];\
					added_1[ 8] <= conv2_bias_array[3];\
					added_1[ 9] <= conv2_bias_array[3];\
					added_1[10] <= conv2_bias_array[3];\
					added_1[11] <= conv2_bias_array[3];\
					added_1[12] <= conv2_bias_array[3];\
					added_1[13] <= conv2_bias_array[3];\
					added_1[14] <= conv2_bias_array[3];\
					added_1[15] <= conv2_bias_array[3];\
					added_1[16] <= conv2_bias_array[3];\
					added_1[17] <= conv2_bias_array[3];\
					added_1[18] <= conv2_bias_array[3];\
					added_1[19] <= conv2_bias_array[3];\
					added_1[20] <= conv2_bias_array[3];\
					added_1[21] <= conv2_bias_array[3];\
					added_1[22] <= conv2_bias_array[3];\
					added_1[23] <= conv2_bias_array[3];\
					added_1[24] <= conv2_bias_array[3];\
					added_1[25] <= conv2_bias_array[3];\
					added_1[26] <= conv2_bias_array[3];\
					added_1[27] <= conv2_bias_array[3];\
					added_1[28] <= conv2_bias_array[3];\
					added_1[29] <= conv2_bias_array[3];\
					added_1[30] <= conv2_bias_array[3];\
					added_1[31] <= conv2_bias_array[3];\
					added_1[32] <= conv2_bias_array[3];\
					added_1[33] <= conv2_bias_array[3];\
					added_1[34] <= conv2_bias_array[3];\
					added_1[35] <= conv2_bias_array[3];\
					added_1[36] <= conv2_bias_array[3];\
					added_1[37] <= conv2_bias_array[3];\
					added_1[38] <= conv2_bias_array[3];\
					added_1[39] <= conv2_bias_array[3];\
					added_1[40] <= conv2_bias_array[3];\
					added_1[41] <= conv2_bias_array[3];\
					added_1[42] <= conv2_bias_array[3];\
					added_1[43] <= conv2_bias_array[3];\
					added_1[44] <= conv2_bias_array[3];\
					added_1[45] <= conv2_bias_array[3];\
					added_1[46] <= conv2_bias_array[3];\
					added_1[47] <= conv2_bias_array[3];\
					added_1[48] <= conv2_bias_array[3];\
					added_1[49] <= conv2_bias_array[3];\
					added_1[50] <= conv2_bias_array[3];\
					added_1[51] <= conv2_bias_array[3];\
					added_1[52] <= conv2_bias_array[3];\
					added_1[53] <= conv2_bias_array[3];\
					added_1[54] <= conv2_bias_array[3];\
					added_1[55] <= conv2_bias_array[3];\
					added_1[56] <= conv2_bias_array[3];\
					added_1[57] <= conv2_bias_array[3];\
					added_1[58] <= conv2_bias_array[3];\
					added_1[59] <= conv2_bias_array[3];\
					added_1[60] <= conv2_bias_array[3];\
					added_1[61] <= conv2_bias_array[3];\
					added_1[62] <= conv2_bias_array[3];\
					added_1[63] <= conv2_bias_array[3];\
					added_1[64] <= conv2_bias_array[3];\
					added_1[65] <= conv2_bias_array[3];\
					added_1[66] <= conv2_bias_array[3];\
					added_1[67] <= conv2_bias_array[3];\
					added_1[68] <= conv2_bias_array[3];\
					added_1[69] <= conv2_bias_array[3];\
					added_1[70] <= conv2_bias_array[3];\
					added_1[71] <= conv2_bias_array[3];\
					added_1[72] <= conv2_bias_array[3];\
					added_1[73] <= conv2_bias_array[3];\
					added_1[74] <= conv2_bias_array[3];\
					added_1[75] <= conv2_bias_array[3];\
					added_1[76] <= conv2_bias_array[3];\
					added_1[77] <= conv2_bias_array[3];\
					added_1[78] <= conv2_bias_array[3];\
					added_1[79] <= conv2_bias_array[3];\
					added_1[80] <= conv2_bias_array[3];\
					added_1[81] <= conv2_bias_array[3];\
					added_1[82] <= conv2_bias_array[3];\
					added_1[83] <= conv2_bias_array[3];\
					added_1[84] <= conv2_bias_array[3];\
					added_1[85] <= conv2_bias_array[3];\
					added_1[86] <= conv2_bias_array[3];\
					added_1[87] <= conv2_bias_array[3];\
					added_1[88] <= conv2_bias_array[3];\
					added_1[89] <= conv2_bias_array[3];\
					added_1[90] <= conv2_bias_array[3];\
					added_1[91] <= conv2_bias_array[3];\
					added_1[92] <= conv2_bias_array[3];\
					added_1[93] <= conv2_bias_array[3];\
					added_1[94] <= conv2_bias_array[3];\
					added_1[95] <= conv2_bias_array[3];\
					added_1[96] <= conv2_bias_array[3];\
					added_1[97] <= conv2_bias_array[3];\
					added_1[98] <= conv2_bias_array[3];\
					added_1[99] <= conv2_bias_array[3];\
				end\
				else begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
				end\
			end\
            CONV2_5_1:begin\
				if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[ 0] <= conv2_bias_array[4];\
					added_1[ 1] <= conv2_bias_array[4];\
					added_1[ 2] <= conv2_bias_array[4];\
					added_1[ 3] <= conv2_bias_array[4];\
					added_1[ 4] <= conv2_bias_array[4];\
					added_1[ 5] <= conv2_bias_array[4];\
					added_1[ 6] <= conv2_bias_array[4];\
					added_1[ 7] <= conv2_bias_array[4];\
					added_1[ 8] <= conv2_bias_array[4];\
					added_1[ 9] <= conv2_bias_array[4];\
					added_1[10] <= conv2_bias_array[4];\
					added_1[11] <= conv2_bias_array[4];\
					added_1[12] <= conv2_bias_array[4];\
					added_1[13] <= conv2_bias_array[4];\
					added_1[14] <= conv2_bias_array[4];\
					added_1[15] <= conv2_bias_array[4];\
					added_1[16] <= conv2_bias_array[4];\
					added_1[17] <= conv2_bias_array[4];\
					added_1[18] <= conv2_bias_array[4];\
					added_1[19] <= conv2_bias_array[4];\
					added_1[20] <= conv2_bias_array[4];\
					added_1[21] <= conv2_bias_array[4];\
					added_1[22] <= conv2_bias_array[4];\
					added_1[23] <= conv2_bias_array[4];\
					added_1[24] <= conv2_bias_array[4];\
					added_1[25] <= conv2_bias_array[4];\
					added_1[26] <= conv2_bias_array[4];\
					added_1[27] <= conv2_bias_array[4];\
					added_1[28] <= conv2_bias_array[4];\
					added_1[29] <= conv2_bias_array[4];\
					added_1[30] <= conv2_bias_array[4];\
					added_1[31] <= conv2_bias_array[4];\
					added_1[32] <= conv2_bias_array[4];\
					added_1[33] <= conv2_bias_array[4];\
					added_1[34] <= conv2_bias_array[4];\
					added_1[35] <= conv2_bias_array[4];\
					added_1[36] <= conv2_bias_array[4];\
					added_1[37] <= conv2_bias_array[4];\
					added_1[38] <= conv2_bias_array[4];\
					added_1[39] <= conv2_bias_array[4];\
					added_1[40] <= conv2_bias_array[4];\
					added_1[41] <= conv2_bias_array[4];\
					added_1[42] <= conv2_bias_array[4];\
					added_1[43] <= conv2_bias_array[4];\
					added_1[44] <= conv2_bias_array[4];\
					added_1[45] <= conv2_bias_array[4];\
					added_1[46] <= conv2_bias_array[4];\
					added_1[47] <= conv2_bias_array[4];\
					added_1[48] <= conv2_bias_array[4];\
					added_1[49] <= conv2_bias_array[4];\
					added_1[50] <= conv2_bias_array[4];\
					added_1[51] <= conv2_bias_array[4];\
					added_1[52] <= conv2_bias_array[4];\
					added_1[53] <= conv2_bias_array[4];\
					added_1[54] <= conv2_bias_array[4];\
					added_1[55] <= conv2_bias_array[4];\
					added_1[56] <= conv2_bias_array[4];\
					added_1[57] <= conv2_bias_array[4];\
					added_1[58] <= conv2_bias_array[4];\
					added_1[59] <= conv2_bias_array[4];\
					added_1[60] <= conv2_bias_array[4];\
					added_1[61] <= conv2_bias_array[4];\
					added_1[62] <= conv2_bias_array[4];\
					added_1[63] <= conv2_bias_array[4];\
					added_1[64] <= conv2_bias_array[4];\
					added_1[65] <= conv2_bias_array[4];\
					added_1[66] <= conv2_bias_array[4];\
					added_1[67] <= conv2_bias_array[4];\
					added_1[68] <= conv2_bias_array[4];\
					added_1[69] <= conv2_bias_array[4];\
					added_1[70] <= conv2_bias_array[4];\
					added_1[71] <= conv2_bias_array[4];\
					added_1[72] <= conv2_bias_array[4];\
					added_1[73] <= conv2_bias_array[4];\
					added_1[74] <= conv2_bias_array[4];\
					added_1[75] <= conv2_bias_array[4];\
					added_1[76] <= conv2_bias_array[4];\
					added_1[77] <= conv2_bias_array[4];\
					added_1[78] <= conv2_bias_array[4];\
					added_1[79] <= conv2_bias_array[4];\
					added_1[80] <= conv2_bias_array[4];\
					added_1[81] <= conv2_bias_array[4];\
					added_1[82] <= conv2_bias_array[4];\
					added_1[83] <= conv2_bias_array[4];\
					added_1[84] <= conv2_bias_array[4];\
					added_1[85] <= conv2_bias_array[4];\
					added_1[86] <= conv2_bias_array[4];\
					added_1[87] <= conv2_bias_array[4];\
					added_1[88] <= conv2_bias_array[4];\
					added_1[89] <= conv2_bias_array[4];\
					added_1[90] <= conv2_bias_array[4];\
					added_1[91] <= conv2_bias_array[4];\
					added_1[92] <= conv2_bias_array[4];\
					added_1[93] <= conv2_bias_array[4];\
					added_1[94] <= conv2_bias_array[4];\
					added_1[95] <= conv2_bias_array[4];\
					added_1[96] <= conv2_bias_array[4];\
					added_1[97] <= conv2_bias_array[4];\
					added_1[98] <= conv2_bias_array[4];\
					added_1[99] <= conv2_bias_array[4];\
				end\
				else begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
				end\
			end\
            CONV2_6_1:begin\
				if((cnt1==8'd0)&(cnt2==8'd0)) begin\
					added_1[ 0] <= conv2_bias_array[5];\
					added_1[ 1] <= conv2_bias_array[5];\
					added_1[ 2] <= conv2_bias_array[5];\
					added_1[ 3] <= conv2_bias_array[5];\
					added_1[ 4] <= conv2_bias_array[5];\
					added_1[ 5] <= conv2_bias_array[5];\
					added_1[ 6] <= conv2_bias_array[5];\
					added_1[ 7] <= conv2_bias_array[5];\
					added_1[ 8] <= conv2_bias_array[5];\
					added_1[ 9] <= conv2_bias_array[5];\
					added_1[10] <= conv2_bias_array[5];\
					added_1[11] <= conv2_bias_array[5];\
					added_1[12] <= conv2_bias_array[5];\
					added_1[13] <= conv2_bias_array[5];\
					added_1[14] <= conv2_bias_array[5];\
					added_1[15] <= conv2_bias_array[5];\
					added_1[16] <= conv2_bias_array[5];\
					added_1[17] <= conv2_bias_array[5];\
					added_1[18] <= conv2_bias_array[5];\
					added_1[19] <= conv2_bias_array[5];\
					added_1[20] <= conv2_bias_array[5];\
					added_1[21] <= conv2_bias_array[5];\
					added_1[22] <= conv2_bias_array[5];\
					added_1[23] <= conv2_bias_array[5];\
					added_1[24] <= conv2_bias_array[5];\
					added_1[25] <= conv2_bias_array[5];\
					added_1[26] <= conv2_bias_array[5];\
					added_1[27] <= conv2_bias_array[5];\
					added_1[28] <= conv2_bias_array[5];\
					added_1[29] <= conv2_bias_array[5];\
					added_1[30] <= conv2_bias_array[5];\
					added_1[31] <= conv2_bias_array[5];\
					added_1[32] <= conv2_bias_array[5];\
					added_1[33] <= conv2_bias_array[5];\
					added_1[34] <= conv2_bias_array[5];\
					added_1[35] <= conv2_bias_array[5];\
					added_1[36] <= conv2_bias_array[5];\
					added_1[37] <= conv2_bias_array[5];\
					added_1[38] <= conv2_bias_array[5];\
					added_1[39] <= conv2_bias_array[5];\
					added_1[40] <= conv2_bias_array[5];\
					added_1[41] <= conv2_bias_array[5];\
					added_1[42] <= conv2_bias_array[5];\
					added_1[43] <= conv2_bias_array[5];\
					added_1[44] <= conv2_bias_array[5];\
					added_1[45] <= conv2_bias_array[5];\
					added_1[46] <= conv2_bias_array[5];\
					added_1[47] <= conv2_bias_array[5];\
					added_1[48] <= conv2_bias_array[5];\
					added_1[49] <= conv2_bias_array[5];\
					added_1[50] <= conv2_bias_array[5];\
					added_1[51] <= conv2_bias_array[5];\
					added_1[52] <= conv2_bias_array[5];\
					added_1[53] <= conv2_bias_array[5];\
					added_1[54] <= conv2_bias_array[5];\
					added_1[55] <= conv2_bias_array[5];\
					added_1[56] <= conv2_bias_array[5];\
					added_1[57] <= conv2_bias_array[5];\
					added_1[58] <= conv2_bias_array[5];\
					added_1[59] <= conv2_bias_array[5];\
					added_1[60] <= conv2_bias_array[5];\
					added_1[61] <= conv2_bias_array[5];\
					added_1[62] <= conv2_bias_array[5];\
					added_1[63] <= conv2_bias_array[5];\
					added_1[64] <= conv2_bias_array[5];\
					added_1[65] <= conv2_bias_array[5];\
					added_1[66] <= conv2_bias_array[5];\
					added_1[67] <= conv2_bias_array[5];\
					added_1[68] <= conv2_bias_array[5];\
					added_1[69] <= conv2_bias_array[5];\
					added_1[70] <= conv2_bias_array[5];\
					added_1[71] <= conv2_bias_array[5];\
					added_1[72] <= conv2_bias_array[5];\
					added_1[73] <= conv2_bias_array[5];\
					added_1[74] <= conv2_bias_array[5];\
					added_1[75] <= conv2_bias_array[5];\
					added_1[76] <= conv2_bias_array[5];\
					added_1[77] <= conv2_bias_array[5];\
					added_1[78] <= conv2_bias_array[5];\
					added_1[79] <= conv2_bias_array[5];\
					added_1[80] <= conv2_bias_array[5];\
					added_1[81] <= conv2_bias_array[5];\
					added_1[82] <= conv2_bias_array[5];\
					added_1[83] <= conv2_bias_array[5];\
					added_1[84] <= conv2_bias_array[5];\
					added_1[85] <= conv2_bias_array[5];\
					added_1[86] <= conv2_bias_array[5];\
					added_1[87] <= conv2_bias_array[5];\
					added_1[88] <= conv2_bias_array[5];\
					added_1[89] <= conv2_bias_array[5];\
					added_1[90] <= conv2_bias_array[5];\
					added_1[91] <= conv2_bias_array[5];\
					added_1[92] <= conv2_bias_array[5];\
					added_1[93] <= conv2_bias_array[5];\
					added_1[94] <= conv2_bias_array[5];\
					added_1[95] <= conv2_bias_array[5];\
					added_1[96] <= conv2_bias_array[5];\
					added_1[97] <= conv2_bias_array[5];\
					added_1[98] <= conv2_bias_array[5];\
					added_1[99] <= conv2_bias_array[5];\
				end\
				else begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
				end\
			end\
            CONV2_1_2,CONV2_1_3,CONV2_1_4,CONV2_1_5,\
			CONV2_2_2,CONV2_2_3,CONV2_2_4,CONV2_2_5,\
			CONV2_3_2,CONV2_3_3,CONV2_3_4,CONV2_3_5,\
			CONV2_4_2,CONV2_4_3,CONV2_4_4,CONV2_4_5,\
			CONV2_5_2,CONV2_5_3,CONV2_5_4,CONV2_5_5,\
			CONV2_6_2,CONV2_6_3,CONV2_6_4,CONV2_6_5:begin\
				added_1[0] <= product_result[0];\
				added_1[1] <= product_result[1];\
				added_1[2] <= product_result[2];\
				added_1[3] <= product_result[3];\
				added_1[4] <= product_result[4];\
				added_1[5] <= product_result[5];\
				added_1[6] <= product_result[6];\
				added_1[7] <= product_result[7];\
				added_1[8] <= product_result[8];\
				added_1[9] <= product_result[9];\
				added_1[10] <= product_result[10];\
				added_1[11] <= product_result[11];\
				added_1[12] <= product_result[12];\
				added_1[13] <= product_result[13];\
				added_1[14] <= product_result[14];\
				added_1[15] <= product_result[15];\
				added_1[16] <= product_result[16];\
				added_1[17] <= product_result[17];\
				added_1[18] <= product_result[18];\
				added_1[19] <= product_result[19];\
				added_1[20] <= product_result[20];\
				added_1[21] <= product_result[21];\
				added_1[22] <= product_result[22];\
				added_1[23] <= product_result[23];\
				added_1[24] <= product_result[24];\
				added_1[25] <= product_result[25];\
				added_1[26] <= product_result[26];\
				added_1[27] <= product_result[27];\
				added_1[28] <= product_result[28];\
				added_1[29] <= product_result[29];\
				added_1[30] <= product_result[30];\
				added_1[31] <= product_result[31];\
				added_1[32] <= product_result[32];\
				added_1[33] <= product_result[33];\
				added_1[34] <= product_result[34];\
				added_1[35] <= product_result[35];\
				added_1[36] <= product_result[36];\
				added_1[37] <= product_result[37];\
				added_1[38] <= product_result[38];\
				added_1[39] <= product_result[39];\
				added_1[40] <= product_result[40];\
				added_1[41] <= product_result[41];\
				added_1[42] <= product_result[42];\
				added_1[43] <= product_result[43];\
				added_1[44] <= product_result[44];\
				added_1[45] <= product_result[45];\
				added_1[46] <= product_result[46];\
				added_1[47] <= product_result[47];\
				added_1[48] <= product_result[48];\
				added_1[49] <= product_result[49];\
				added_1[50] <= product_result[50];\
				added_1[51] <= product_result[51];\
				added_1[52] <= product_result[52];\
				added_1[53] <= product_result[53];\
				added_1[54] <= product_result[54];\
				added_1[55] <= product_result[55];\
				added_1[56] <= product_result[56];\
				added_1[57] <= product_result[57];\
				added_1[58] <= product_result[58];\
				added_1[59] <= product_result[59];\
				added_1[60] <= product_result[60];\
				added_1[61] <= product_result[61];\
				added_1[62] <= product_result[62];\
				added_1[63] <= product_result[63];\
				added_1[64] <= product_result[64];\
				added_1[65] <= product_result[65];\
				added_1[66] <= product_result[66];\
				added_1[67] <= product_result[67];\
				added_1[68] <= product_result[68];\
				added_1[69] <= product_result[69];\
				added_1[70] <= product_result[70];\
				added_1[71] <= product_result[71];\
				added_1[72] <= product_result[72];\
				added_1[73] <= product_result[73];\
				added_1[74] <= product_result[74];\
				added_1[75] <= product_result[75];\
				added_1[76] <= product_result[76];\
				added_1[77] <= product_result[77];\
				added_1[78] <= product_result[78];\
				added_1[79] <= product_result[79];\
				added_1[80] <= product_result[80];\
				added_1[81] <= product_result[81];\
				added_1[82] <= product_result[82];\
				added_1[83] <= product_result[83];\
				added_1[84] <= product_result[84];\
				added_1[85] <= product_result[85];\
				added_1[86] <= product_result[86];\
				added_1[87] <= product_result[87];\
				added_1[88] <= product_result[88];\
				added_1[89] <= product_result[89];\
				added_1[90] <= product_result[90];\
				added_1[91] <= product_result[91];\
				added_1[92] <= product_result[92];\
				added_1[93] <= product_result[93];\
				added_1[94] <= product_result[94];\
				added_1[95] <= product_result[95];\
				added_1[96] <= product_result[96];\
				added_1[97] <= product_result[97];\
				added_1[98] <= product_result[98];\
				added_1[99] <= product_result[99];\
				added_2[0] <= add_result[0];\
				added_2[1] <= add_result[1];\
				added_2[2] <= add_result[2];\
				added_2[3] <= add_result[3];\
				added_2[4] <= add_result[4];\
				added_2[5] <= add_result[5];\
				added_2[6] <= add_result[6];\
				added_2[7] <= add_result[7];\
				added_2[8] <= add_result[8];\
				added_2[9] <= add_result[9];\
				added_2[10] <= add_result[10];\
				added_2[11] <= add_result[11];\
				added_2[12] <= add_result[12];\
				added_2[13] <= add_result[13];\
				added_2[14] <= add_result[14];\
				added_2[15] <= add_result[15];\
				added_2[16] <= add_result[16];\
				added_2[17] <= add_result[17];\
				added_2[18] <= add_result[18];\
				added_2[19] <= add_result[19];\
				added_2[20] <= add_result[20];\
				added_2[21] <= add_result[21];\
				added_2[22] <= add_result[22];\
				added_2[23] <= add_result[23];\
				added_2[24] <= add_result[24];\
				added_2[25] <= add_result[25];\
				added_2[26] <= add_result[26];\
				added_2[27] <= add_result[27];\
				added_2[28] <= add_result[28];\
				added_2[29] <= add_result[29];\
				added_2[30] <= add_result[30];\
				added_2[31] <= add_result[31];\
				added_2[32] <= add_result[32];\
				added_2[33] <= add_result[33];\
				added_2[34] <= add_result[34];\
				added_2[35] <= add_result[35];\
				added_2[36] <= add_result[36];\
				added_2[37] <= add_result[37];\
				added_2[38] <= add_result[38];\
				added_2[39] <= add_result[39];\
				added_2[40] <= add_result[40];\
				added_2[41] <= add_result[41];\
				added_2[42] <= add_result[42];\
				added_2[43] <= add_result[43];\
				added_2[44] <= add_result[44];\
				added_2[45] <= add_result[45];\
				added_2[46] <= add_result[46];\
				added_2[47] <= add_result[47];\
				added_2[48] <= add_result[48];\
				added_2[49] <= add_result[49];\
				added_2[50] <= add_result[50];\
				added_2[51] <= add_result[51];\
				added_2[52] <= add_result[52];\
				added_2[53] <= add_result[53];\
				added_2[54] <= add_result[54];\
				added_2[55] <= add_result[55];\
				added_2[56] <= add_result[56];\
				added_2[57] <= add_result[57];\
				added_2[58] <= add_result[58];\
				added_2[59] <= add_result[59];\
				added_2[60] <= add_result[60];\
				added_2[61] <= add_result[61];\
				added_2[62] <= add_result[62];\
				added_2[63] <= add_result[63];\
				added_2[64] <= add_result[64];\
				added_2[65] <= add_result[65];\
				added_2[66] <= add_result[66];\
				added_2[67] <= add_result[67];\
				added_2[68] <= add_result[68];\
				added_2[69] <= add_result[69];\
				added_2[70] <= add_result[70];\
				added_2[71] <= add_result[71];\
				added_2[72] <= add_result[72];\
				added_2[73] <= add_result[73];\
				added_2[74] <= add_result[74];\
				added_2[75] <= add_result[75];\
				added_2[76] <= add_result[76];\
				added_2[77] <= add_result[77];\
				added_2[78] <= add_result[78];\
				added_2[79] <= add_result[79];\
				added_2[80] <= add_result[80];\
				added_2[81] <= add_result[81];\
				added_2[82] <= add_result[82];\
				added_2[83] <= add_result[83];\
				added_2[84] <= add_result[84];\
				added_2[85] <= add_result[85];\
				added_2[86] <= add_result[86];\
				added_2[87] <= add_result[87];\
				added_2[88] <= add_result[88];\
				added_2[89] <= add_result[89];\
				added_2[90] <= add_result[90];\
				added_2[91] <= add_result[91];\
				added_2[92] <= add_result[92];\
				added_2[93] <= add_result[93];\
				added_2[94] <= add_result[94];\
				added_2[95] <= add_result[95];\
				added_2[96] <= add_result[96];\
				added_2[97] <= add_result[97];\
				added_2[98] <= add_result[98];\
				added_2[99] <= add_result[99];\
			end\
            CONV2_1_6,CONV2_2_6,CONV2_3_6,CONV2_4_6,CONV2_5_6,CONV2_6_6:begin\
				if(cnt2<8'd6)begin\
					added_1[0] <= product_result[0];\
					added_1[1] <= product_result[1];\
					added_1[2] <= product_result[2];\
					added_1[3] <= product_result[3];\
					added_1[4] <= product_result[4];\
					added_1[5] <= product_result[5];\
					added_1[6] <= product_result[6];\
					added_1[7] <= product_result[7];\
					added_1[8] <= product_result[8];\
					added_1[9] <= product_result[9];\
					added_1[10] <= product_result[10];\
					added_1[11] <= product_result[11];\
					added_1[12] <= product_result[12];\
					added_1[13] <= product_result[13];\
					added_1[14] <= product_result[14];\
					added_1[15] <= product_result[15];\
					added_1[16] <= product_result[16];\
					added_1[17] <= product_result[17];\
					added_1[18] <= product_result[18];\
					added_1[19] <= product_result[19];\
					added_1[20] <= product_result[20];\
					added_1[21] <= product_result[21];\
					added_1[22] <= product_result[22];\
					added_1[23] <= product_result[23];\
					added_1[24] <= product_result[24];\
					added_1[25] <= product_result[25];\
					added_1[26] <= product_result[26];\
					added_1[27] <= product_result[27];\
					added_1[28] <= product_result[28];\
					added_1[29] <= product_result[29];\
					added_1[30] <= product_result[30];\
					added_1[31] <= product_result[31];\
					added_1[32] <= product_result[32];\
					added_1[33] <= product_result[33];\
					added_1[34] <= product_result[34];\
					added_1[35] <= product_result[35];\
					added_1[36] <= product_result[36];\
					added_1[37] <= product_result[37];\
					added_1[38] <= product_result[38];\
					added_1[39] <= product_result[39];\
					added_1[40] <= product_result[40];\
					added_1[41] <= product_result[41];\
					added_1[42] <= product_result[42];\
					added_1[43] <= product_result[43];\
					added_1[44] <= product_result[44];\
					added_1[45] <= product_result[45];\
					added_1[46] <= product_result[46];\
					added_1[47] <= product_result[47];\
					added_1[48] <= product_result[48];\
					added_1[49] <= product_result[49];\
					added_1[50] <= product_result[50];\
					added_1[51] <= product_result[51];\
					added_1[52] <= product_result[52];\
					added_1[53] <= product_result[53];\
					added_1[54] <= product_result[54];\
					added_1[55] <= product_result[55];\
					added_1[56] <= product_result[56];\
					added_1[57] <= product_result[57];\
					added_1[58] <= product_result[58];\
					added_1[59] <= product_result[59];\
					added_1[60] <= product_result[60];\
					added_1[61] <= product_result[61];\
					added_1[62] <= product_result[62];\
					added_1[63] <= product_result[63];\
					added_1[64] <= product_result[64];\
					added_1[65] <= product_result[65];\
					added_1[66] <= product_result[66];\
					added_1[67] <= product_result[67];\
					added_1[68] <= product_result[68];\
					added_1[69] <= product_result[69];\
					added_1[70] <= product_result[70];\
					added_1[71] <= product_result[71];\
					added_1[72] <= product_result[72];\
					added_1[73] <= product_result[73];\
					added_1[74] <= product_result[74];\
					added_1[75] <= product_result[75];\
					added_1[76] <= product_result[76];\
					added_1[77] <= product_result[77];\
					added_1[78] <= product_result[78];\
					added_1[79] <= product_result[79];\
					added_1[80] <= product_result[80];\
					added_1[81] <= product_result[81];\
					added_1[82] <= product_result[82];\
					added_1[83] <= product_result[83];\
					added_1[84] <= product_result[84];\
					added_1[85] <= product_result[85];\
					added_1[86] <= product_result[86];\
					added_1[87] <= product_result[87];\
					added_1[88] <= product_result[88];\
					added_1[89] <= product_result[89];\
					added_1[90] <= product_result[90];\
					added_1[91] <= product_result[91];\
					added_1[92] <= product_result[92];\
					added_1[93] <= product_result[93];\
					added_1[94] <= product_result[94];\
					added_1[95] <= product_result[95];\
					added_1[96] <= product_result[96];\
					added_1[97] <= product_result[97];\
					added_1[98] <= product_result[98];\
					added_1[99] <= product_result[99];\
					added_2[0] <= add_result[0];\
					added_2[1] <= add_result[1];\
					added_2[2] <= add_result[2];\
					added_2[3] <= add_result[3];\
					added_2[4] <= add_result[4];\
					added_2[5] <= add_result[5];\
					added_2[6] <= add_result[6];\
					added_2[7] <= add_result[7];\
					added_2[8] <= add_result[8];\
					added_2[9] <= add_result[9];\
					added_2[10] <= add_result[10];\
					added_2[11] <= add_result[11];\
					added_2[12] <= add_result[12];\
					added_2[13] <= add_result[13];\
					added_2[14] <= add_result[14];\
					added_2[15] <= add_result[15];\
					added_2[16] <= add_result[16];\
					added_2[17] <= add_result[17];\
					added_2[18] <= add_result[18];\
					added_2[19] <= add_result[19];\
					added_2[20] <= add_result[20];\
					added_2[21] <= add_result[21];\
					added_2[22] <= add_result[22];\
					added_2[23] <= add_result[23];\
					added_2[24] <= add_result[24];\
					added_2[25] <= add_result[25];\
					added_2[26] <= add_result[26];\
					added_2[27] <= add_result[27];\
					added_2[28] <= add_result[28];\
					added_2[29] <= add_result[29];\
					added_2[30] <= add_result[30];\
					added_2[31] <= add_result[31];\
					added_2[32] <= add_result[32];\
					added_2[33] <= add_result[33];\
					added_2[34] <= add_result[34];\
					added_2[35] <= add_result[35];\
					added_2[36] <= add_result[36];\
					added_2[37] <= add_result[37];\
					added_2[38] <= add_result[38];\
					added_2[39] <= add_result[39];\
					added_2[40] <= add_result[40];\
					added_2[41] <= add_result[41];\
					added_2[42] <= add_result[42];\
					added_2[43] <= add_result[43];\
					added_2[44] <= add_result[44];\
					added_2[45] <= add_result[45];\
					added_2[46] <= add_result[46];\
					added_2[47] <= add_result[47];\
					added_2[48] <= add_result[48];\
					added_2[49] <= add_result[49];\
					added_2[50] <= add_result[50];\
					added_2[51] <= add_result[51];\
					added_2[52] <= add_result[52];\
					added_2[53] <= add_result[53];\
					added_2[54] <= add_result[54];\
					added_2[55] <= add_result[55];\
					added_2[56] <= add_result[56];\
					added_2[57] <= add_result[57];\
					added_2[58] <= add_result[58];\
					added_2[59] <= add_result[59];\
					added_2[60] <= add_result[60];\
					added_2[61] <= add_result[61];\
					added_2[62] <= add_result[62];\
					added_2[63] <= add_result[63];\
					added_2[64] <= add_result[64];\
					added_2[65] <= add_result[65];\
					added_2[66] <= add_result[66];\
					added_2[67] <= add_result[67];\
					added_2[68] <= add_result[68];\
					added_2[69] <= add_result[69];\
					added_2[70] <= add_result[70];\
					added_2[71] <= add_result[71];\
					added_2[72] <= add_result[72];\
					added_2[73] <= add_result[73];\
					added_2[74] <= add_result[74];\
					added_2[75] <= add_result[75];\
					added_2[76] <= add_result[76];\
					added_2[77] <= add_result[77];\
					added_2[78] <= add_result[78];\
					added_2[79] <= add_result[79];\
					added_2[80] <= add_result[80];\
					added_2[81] <= add_result[81];\
					added_2[82] <= add_result[82];\
					added_2[83] <= add_result[83];\
					added_2[84] <= add_result[84];\
					added_2[85] <= add_result[85];\
					added_2[86] <= add_result[86];\
					added_2[87] <= add_result[87];\
					added_2[88] <= add_result[88];\
					added_2[89] <= add_result[89];\
					added_2[90] <= add_result[90];\
					added_2[91] <= add_result[91];\
					added_2[92] <= add_result[92];\
					added_2[93] <= add_result[93];\
					added_2[94] <= add_result[94];\
					added_2[95] <= add_result[95];\
					added_2[96] <= add_result[96];\
					added_2[97] <= add_result[97];\
					added_2[98] <= add_result[98];\
					added_2[99] <= add_result[99];\
				end\
				else begin\
                    added_2[0] <= 18'd0;\
                    added_2[1] <= 18'd0;\
                    added_2[2] <= 18'd0;\
                    added_2[3] <= 18'd0;\
                    added_2[4] <= 18'd0;\
                    added_2[5] <= 18'd0;\
                    added_2[6] <= 18'd0;\
                    added_2[7] <= 18'd0;\
                    added_2[8] <= 18'd0;\
                    added_2[9] <= 18'd0;\
                    added_2[10] <= 18'd0;\
                    added_2[11] <= 18'd0;\
                    added_2[12] <= 18'd0;\
                    added_2[13] <= 18'd0;\
                    added_2[14] <= 18'd0;\
                    added_2[15] <= 18'd0;\
                    added_2[16] <= 18'd0;\
                    added_2[17] <= 18'd0;\
                    added_2[18] <= 18'd0;\
                    added_2[19] <= 18'd0;\
                    added_2[20] <= 18'd0;\
                    added_2[21] <= 18'd0;\
                    added_2[22] <= 18'd0;\
                    added_2[23] <= 18'd0;\
                    added_2[24] <= 18'd0;\
                    added_2[25] <= 18'd0;\
                    added_2[26] <= 18'd0;\
                    added_2[27] <= 18'd0;\
                    added_2[28] <= 18'd0;\
                    added_2[29] <= 18'd0;\
                    added_2[30] <= 18'd0;\
                    added_2[31] <= 18'd0;\
                    added_2[32] <= 18'd0;\
                    added_2[33] <= 18'd0;\
                    added_2[34] <= 18'd0;\
                    added_2[35] <= 18'd0;\
                    added_2[36] <= 18'd0;\
                    added_2[37] <= 18'd0;\
                    added_2[38] <= 18'd0;\
                    added_2[39] <= 18'd0;\
                    added_2[40] <= 18'd0;\
                    added_2[41] <= 18'd0;\
                    added_2[42] <= 18'd0;\
                    added_2[43] <= 18'd0;\
                    added_2[44] <= 18'd0;\
                    added_2[45] <= 18'd0;\
                    added_2[46] <= 18'd0;\
                    added_2[47] <= 18'd0;\
                    added_2[48] <= 18'd0;\
                    added_2[49] <= 18'd0;\
                    added_2[50] <= 18'd0;\
                    added_2[51] <= 18'd0;\
                    added_2[52] <= 18'd0;\
                    added_2[53] <= 18'd0;\
                    added_2[54] <= 18'd0;\
                    added_2[55] <= 18'd0;\
                    added_2[56] <= 18'd0;\
                    added_2[57] <= 18'd0;\
                    added_2[58] <= 18'd0;\
                    added_2[59] <= 18'd0;\
                    added_2[60] <= 18'd0;\
                    added_2[61] <= 18'd0;\
                    added_2[62] <= 18'd0;\
                    added_2[63] <= 18'd0;\
                    added_2[64] <= 18'd0;\
                    added_2[65] <= 18'd0;\
                    added_2[66] <= 18'd0;\
                    added_2[67] <= 18'd0;\
                    added_2[68] <= 18'd0;\
                    added_2[69] <= 18'd0;\
                    added_2[70] <= 18'd0;\
                    added_2[71] <= 18'd0;\
                    added_2[72] <= 18'd0;\
                    added_2[73] <= 18'd0;\
                    added_2[74] <= 18'd0;\
                    added_2[75] <= 18'd0;\
                    added_2[76] <= 18'd0;\
                    added_2[77] <= 18'd0;\
                    added_2[78] <= 18'd0;\
                    added_2[79] <= 18'd0;\
                    added_2[80] <= 18'd0;\
                    added_2[81] <= 18'd0;\
                    added_2[82] <= 18'd0;\
                    added_2[83] <= 18'd0;\
                    added_2[84] <= 18'd0;\
                    added_2[85] <= 18'd0;\
                    added_2[86] <= 18'd0;\
                    added_2[87] <= 18'd0;\
                    added_2[88] <= 18'd0;\
                    added_2[89] <= 18'd0;\
                    added_2[90] <= 18'd0;\
                    added_2[91] <= 18'd0;\
                    added_2[92] <= 18'd0;\
                    added_2[93] <= 18'd0;\
                    added_2[94] <= 18'd0;\
                    added_2[95] <= 18'd0;\
                    added_2[96] <= 18'd0;\
                    added_2[97] <= 18'd0;\
                    added_2[98] <= 18'd0;\
                    added_2[99] <= 18'd0;\
                end\
			end\
            LINEAR1  :begin\
				if(cnt1==8'd0) begin\
					added_1[100] <= linear1_bias_array[0];\
					added_1[101] <= linear1_bias_array[1];\
					added_1[102] <= linear1_bias_array[2];\
					added_1[103] <= linear1_bias_array[3];\
					added_1[104] <= linear1_bias_array[4];\
					added_1[105] <= linear1_bias_array[5];\
					added_1[106] <= linear1_bias_array[6];\
					added_1[107] <= linear1_bias_array[7];\
					added_1[108] <= linear1_bias_array[8];\
					added_1[109] <= linear1_bias_array[9];\
					added_1[110] <= linear1_bias_array[10];\
					added_1[111] <= linear1_bias_array[11];\
				end\
				else if(cnt1<8'd151) begin\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_1[110] <= product_result[110];\
					added_1[111] <= product_result[111];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
					added_2[110] <= add_result[110];\
					added_2[111] <= add_result[111];\
				end\
				else begin\
					added_1[100] <= 18'd0;\
					added_1[101] <= 18'd0;\
					added_1[102] <= 18'd0;\
					added_1[103] <= 18'd0;\
					added_1[104] <= 18'd0;\
					added_1[105] <= 18'd0;\
					added_1[106] <= 18'd0;\
					added_1[107] <= 18'd0;\
					added_1[108] <= 18'd0;\
					added_1[109] <= 18'd0;\
					added_1[110] <= 18'd0;\
					added_1[111] <= 18'd0;\
					added_2[100] <= 18'd0;\
					added_2[101] <= 18'd0;\
					added_2[102] <= 18'd0;\
					added_2[103] <= 18'd0;\
					added_2[104] <= 18'd0;\
					added_2[105] <= 18'd0;\
					added_2[106] <= 18'd0;\
					added_2[107] <= 18'd0;\
					added_2[108] <= 18'd0;\
					added_2[109] <= 18'd0;\
					added_2[110] <= 18'd0;\
					added_2[111] <= 18'd0;\
				end\
			end\
            LINEAR2  :begin\
				if(cnt2==8'd0)begin\
					added_1[100] <= linear2_bias_array[0];\
					added_1[101] <= linear2_bias_array[1];\
					added_1[102] <= linear2_bias_array[2];\
					added_1[103] <= linear2_bias_array[3];\
					added_1[104] <= linear2_bias_array[4];\
					added_1[105] <= linear2_bias_array[5];\
					added_1[106] <= linear2_bias_array[6];\
					added_1[107] <= linear2_bias_array[7];\
					added_1[108] <= linear2_bias_array[8];\
					added_1[109] <= linear2_bias_array[9];\
				end\
				else if(cnt2<8'd13)begin\
					added_1[100] <= product_result[100];\
					added_1[101] <= product_result[101];\
					added_1[102] <= product_result[102];\
					added_1[103] <= product_result[103];\
					added_1[104] <= product_result[104];\
					added_1[105] <= product_result[105];\
					added_1[106] <= product_result[106];\
					added_1[107] <= product_result[107];\
					added_1[108] <= product_result[108];\
					added_1[109] <= product_result[109];\
					added_2[100] <= add_result[100];\
					added_2[101] <= add_result[101];\
					added_2[102] <= add_result[102];\
					added_2[103] <= add_result[103];\
					added_2[104] <= add_result[104];\
					added_2[105] <= add_result[105];\
					added_2[106] <= add_result[106];\
					added_2[107] <= add_result[107];\
					added_2[108] <= add_result[108];\
					added_2[109] <= add_result[109];\
				end\
				else begin\
					added_1[100] <= 18'd0;\
					added_1[101] <= 18'd0;\
					added_1[102] <= 18'd0;\
					added_1[103] <= 18'd0;\
					added_1[104] <= 18'd0;\
					added_1[105] <= 18'd0;\
					added_1[106] <= 18'd0;\
					added_1[107] <= 18'd0;\
					added_1[108] <= 18'd0;\
					added_1[109] <= 18'd0;\
					added_2[100] <= 18'd0;\
					added_2[101] <= 18'd0;\
					added_2[102] <= 18'd0;\
					added_2[103] <= 18'd0;\
					added_2[104] <= 18'd0;\
					added_2[105] <= 18'd0;\
					added_2[106] <= 18'd0;\
					added_2[107] <= 18'd0;\
					added_2[108] <= 18'd0;\
					added_2[109] <= 18'd0;\
				end\
			end\
			COMPARE  :;\
            COMPLETE :;\
            default: begin\
				added_1[0] <= 18'd0;\
				added_1[1] <= 18'd0;\
				added_1[2] <= 18'd0;\
				added_1[3] <= 18'd0;\
				added_1[4] <= 18'd0;\
				added_1[5] <= 18'd0;\
				added_1[6] <= 18'd0;\
				added_1[7] <= 18'd0;\
				added_1[8] <= 18'd0;\
				added_1[9] <= 18'd0;\
				added_1[10] <= 18'd0;\
				added_1[11] <= 18'd0;\
				added_1[12] <= 18'd0;\
				added_1[13] <= 18'd0;\
				added_1[14] <= 18'd0;\
				added_1[15] <= 18'd0;\
				added_1[16] <= 18'd0;\
				added_1[17] <= 18'd0;\
				added_1[18] <= 18'd0;\
				added_1[19] <= 18'd0;\
				added_1[20] <= 18'd0;\
				added_1[21] <= 18'd0;\
				added_1[22] <= 18'd0;\
				added_1[23] <= 18'd0;\
				added_1[24] <= 18'd0;\
				added_1[25] <= 18'd0;\
				added_1[26] <= 18'd0;\
				added_1[27] <= 18'd0;\
				added_1[28] <= 18'd0;\
				added_1[29] <= 18'd0;\
				added_1[30] <= 18'd0;\
				added_1[31] <= 18'd0;\
				added_1[32] <= 18'd0;\
				added_1[33] <= 18'd0;\
				added_1[34] <= 18'd0;\
				added_1[35] <= 18'd0;\
				added_1[36] <= 18'd0;\
				added_1[37] <= 18'd0;\
				added_1[38] <= 18'd0;\
				added_1[39] <= 18'd0;\
				added_1[40] <= 18'd0;\
				added_1[41] <= 18'd0;\
				added_1[42] <= 18'd0;\
				added_1[43] <= 18'd0;\
				added_1[44] <= 18'd0;\
				added_1[45] <= 18'd0;\
				added_1[46] <= 18'd0;\
				added_1[47] <= 18'd0;\
				added_1[48] <= 18'd0;\
				added_1[49] <= 18'd0;\
				added_1[50] <= 18'd0;\
				added_1[51] <= 18'd0;\
				added_1[52] <= 18'd0;\
				added_1[53] <= 18'd0;\
				added_1[54] <= 18'd0;\
				added_1[55] <= 18'd0;\
				added_1[56] <= 18'd0;\
				added_1[57] <= 18'd0;\
				added_1[58] <= 18'd0;\
				added_1[59] <= 18'd0;\
				added_1[60] <= 18'd0;\
				added_1[61] <= 18'd0;\
				added_1[62] <= 18'd0;\
				added_1[63] <= 18'd0;\
				added_1[64] <= 18'd0;\
				added_1[65] <= 18'd0;\
				added_1[66] <= 18'd0;\
				added_1[67] <= 18'd0;\
				added_1[68] <= 18'd0;\
				added_1[69] <= 18'd0;\
				added_1[70] <= 18'd0;\
				added_1[71] <= 18'd0;\
				added_1[72] <= 18'd0;\
				added_1[73] <= 18'd0;\
				added_1[74] <= 18'd0;\
				added_1[75] <= 18'd0;\
				added_1[76] <= 18'd0;\
				added_1[77] <= 18'd0;\
				added_1[78] <= 18'd0;\
				added_1[79] <= 18'd0;\
				added_1[80] <= 18'd0;\
				added_1[81] <= 18'd0;\
				added_1[82] <= 18'd0;\
				added_1[83] <= 18'd0;\
				added_1[84] <= 18'd0;\
				added_1[85] <= 18'd0;\
				added_1[86] <= 18'd0;\
				added_1[87] <= 18'd0;\
				added_1[88] <= 18'd0;\
				added_1[89] <= 18'd0;\
				added_1[90] <= 18'd0;\
				added_1[91] <= 18'd0;\
				added_1[92] <= 18'd0;\
				added_1[93] <= 18'd0;\
				added_1[94] <= 18'd0;\
				added_1[95] <= 18'd0;\
				added_1[96] <= 18'd0;\
				added_1[97] <= 18'd0;\
				added_1[98] <= 18'd0;\
				added_1[99] <= 18'd0;\
				added_1[100] <= 18'd0;\
				added_1[101] <= 18'd0;\
				added_1[102] <= 18'd0;\
				added_1[103] <= 18'd0;\
				added_1[104] <= 18'd0;\
				added_1[105] <= 18'd0;\
				added_1[106] <= 18'd0;\
				added_1[107] <= 18'd0;\
				added_1[108] <= 18'd0;\
				added_1[109] <= 18'd0;\
				added_1[110] <= 18'd0;\
				added_1[111] <= 18'd0;\
				added_2[0] <= 18'd0;\
				added_2[1] <= 18'd0;\
				added_2[2] <= 18'd0;\
				added_2[3] <= 18'd0;\
				added_2[4] <= 18'd0;\
				added_2[5] <= 18'd0;\
				added_2[6] <= 18'd0;\
				added_2[7] <= 18'd0;\
				added_2[8] <= 18'd0;\
				added_2[9] <= 18'd0;\
				added_2[10] <= 18'd0;\
				added_2[11] <= 18'd0;\
				added_2[12] <= 18'd0;\
				added_2[13] <= 18'd0;\
				added_2[14] <= 18'd0;\
				added_2[15] <= 18'd0;\
				added_2[16] <= 18'd0;\
				added_2[17] <= 18'd0;\
				added_2[18] <= 18'd0;\
				added_2[19] <= 18'd0;\
				added_2[20] <= 18'd0;\
				added_2[21] <= 18'd0;\
				added_2[22] <= 18'd0;\
				added_2[23] <= 18'd0;\
				added_2[24] <= 18'd0;\
				added_2[25] <= 18'd0;\
				added_2[26] <= 18'd0;\
				added_2[27] <= 18'd0;\
				added_2[28] <= 18'd0;\
				added_2[29] <= 18'd0;\
				added_2[30] <= 18'd0;\
				added_2[31] <= 18'd0;\
				added_2[32] <= 18'd0;\
				added_2[33] <= 18'd0;\
				added_2[34] <= 18'd0;\
				added_2[35] <= 18'd0;\
				added_2[36] <= 18'd0;\
				added_2[37] <= 18'd0;\
				added_2[38] <= 18'd0;\
				added_2[39] <= 18'd0;\
				added_2[40] <= 18'd0;\
				added_2[41] <= 18'd0;\
				added_2[42] <= 18'd0;\
				added_2[43] <= 18'd0;\
				added_2[44] <= 18'd0;\
				added_2[45] <= 18'd0;\
				added_2[46] <= 18'd0;\
				added_2[47] <= 18'd0;\
				added_2[48] <= 18'd0;\
				added_2[49] <= 18'd0;\
				added_2[50] <= 18'd0;\
				added_2[51] <= 18'd0;\
				added_2[52] <= 18'd0;\
				added_2[53] <= 18'd0;\
				added_2[54] <= 18'd0;\
				added_2[55] <= 18'd0;\
				added_2[56] <= 18'd0;\
				added_2[57] <= 18'd0;\
				added_2[58] <= 18'd0;\
				added_2[59] <= 18'd0;\
				added_2[60] <= 18'd0;\
				added_2[61] <= 18'd0;\
				added_2[62] <= 18'd0;\
				added_2[63] <= 18'd0;\
				added_2[64] <= 18'd0;\
				added_2[65] <= 18'd0;\
				added_2[66] <= 18'd0;\
				added_2[67] <= 18'd0;\
				added_2[68] <= 18'd0;\
				added_2[69] <= 18'd0;\
				added_2[70] <= 18'd0;\
				added_2[71] <= 18'd0;\
				added_2[72] <= 18'd0;\
				added_2[73] <= 18'd0;\
				added_2[74] <= 18'd0;\
				added_2[75] <= 18'd0;\
				added_2[76] <= 18'd0;\
				added_2[77] <= 18'd0;\
				added_2[78] <= 18'd0;\
				added_2[79] <= 18'd0;\
				added_2[80] <= 18'd0;\
				added_2[81] <= 18'd0;\
				added_2[82] <= 18'd0;\
				added_2[83] <= 18'd0;\
				added_2[84] <= 18'd0;\
				added_2[85] <= 18'd0;\
				added_2[86] <= 18'd0;\
				added_2[87] <= 18'd0;\
				added_2[88] <= 18'd0;\
				added_2[89] <= 18'd0;\
				added_2[90] <= 18'd0;\
				added_2[91] <= 18'd0;\
				added_2[92] <= 18'd0;\
				added_2[93] <= 18'd0;\
				added_2[94] <= 18'd0;\
				added_2[95] <= 18'd0;\
				added_2[96] <= 18'd0;\
				added_2[97] <= 18'd0;\
				added_2[98] <= 18'd0;\
				added_2[99] <= 18'd0;\
				added_2[100] <= 18'd0;\
				added_2[101] <= 18'd0;\
				added_2[102] <= 18'd0;\
				added_2[103] <= 18'd0;\
				added_2[104] <= 18'd0;\
				added_2[105] <= 18'd0;\
				added_2[106] <= 18'd0;\
				added_2[107] <= 18'd0;\
				added_2[108] <= 18'd0;\
				added_2[109] <= 18'd0;\
				added_2[110] <= 18'd0;\
				added_2[111] <= 18'd0;\
			end\
        endcase\
    end\
end