`define CONV1_RESULT \
always@(posedge clk or negedge rst_n) begin\
    if(!rst_n)begin\
		conv1_result[0][0][0] <= 18'd0;\
		conv1_result[0][0][1] <= 18'd0;\
		conv1_result[0][0][2] <= 18'd0;\
		conv1_result[0][0][3] <= 18'd0;\
		conv1_result[0][0][4] <= 18'd0;\
		conv1_result[0][0][5] <= 18'd0;\
		conv1_result[0][0][6] <= 18'd0;\
		conv1_result[0][0][7] <= 18'd0;\
		conv1_result[0][0][8] <= 18'd0;\
		conv1_result[0][0][9] <= 18'd0;\
		conv1_result[0][0][10] <= 18'd0;\
		conv1_result[0][0][11] <= 18'd0;\
		conv1_result[0][0][12] <= 18'd0;\
		conv1_result[0][0][13] <= 18'd0;\
		conv1_result[0][1][0] <= 18'd0;\
		conv1_result[0][1][1] <= 18'd0;\
		conv1_result[0][1][2] <= 18'd0;\
		conv1_result[0][1][3] <= 18'd0;\
		conv1_result[0][1][4] <= 18'd0;\
		conv1_result[0][1][5] <= 18'd0;\
		conv1_result[0][1][6] <= 18'd0;\
		conv1_result[0][1][7] <= 18'd0;\
		conv1_result[0][1][8] <= 18'd0;\
		conv1_result[0][1][9] <= 18'd0;\
		conv1_result[0][1][10] <= 18'd0;\
		conv1_result[0][1][11] <= 18'd0;\
		conv1_result[0][1][12] <= 18'd0;\
		conv1_result[0][1][13] <= 18'd0;\
		conv1_result[0][2][0] <= 18'd0;\
		conv1_result[0][2][1] <= 18'd0;\
		conv1_result[0][2][2] <= 18'd0;\
		conv1_result[0][2][3] <= 18'd0;\
		conv1_result[0][2][4] <= 18'd0;\
		conv1_result[0][2][5] <= 18'd0;\
		conv1_result[0][2][6] <= 18'd0;\
		conv1_result[0][2][7] <= 18'd0;\
		conv1_result[0][2][8] <= 18'd0;\
		conv1_result[0][2][9] <= 18'd0;\
		conv1_result[0][2][10] <= 18'd0;\
		conv1_result[0][2][11] <= 18'd0;\
		conv1_result[0][2][12] <= 18'd0;\
		conv1_result[0][2][13] <= 18'd0;\
		conv1_result[0][3][0] <= 18'd0;\
		conv1_result[0][3][1] <= 18'd0;\
		conv1_result[0][3][2] <= 18'd0;\
		conv1_result[0][3][3] <= 18'd0;\
		conv1_result[0][3][4] <= 18'd0;\
		conv1_result[0][3][5] <= 18'd0;\
		conv1_result[0][3][6] <= 18'd0;\
		conv1_result[0][3][7] <= 18'd0;\
		conv1_result[0][3][8] <= 18'd0;\
		conv1_result[0][3][9] <= 18'd0;\
		conv1_result[0][3][10] <= 18'd0;\
		conv1_result[0][3][11] <= 18'd0;\
		conv1_result[0][3][12] <= 18'd0;\
		conv1_result[0][3][13] <= 18'd0;\
		conv1_result[0][4][0] <= 18'd0;\
		conv1_result[0][4][1] <= 18'd0;\
		conv1_result[0][4][2] <= 18'd0;\
		conv1_result[0][4][3] <= 18'd0;\
		conv1_result[0][4][4] <= 18'd0;\
		conv1_result[0][4][5] <= 18'd0;\
		conv1_result[0][4][6] <= 18'd0;\
		conv1_result[0][4][7] <= 18'd0;\
		conv1_result[0][4][8] <= 18'd0;\
		conv1_result[0][4][9] <= 18'd0;\
		conv1_result[0][4][10] <= 18'd0;\
		conv1_result[0][4][11] <= 18'd0;\
		conv1_result[0][4][12] <= 18'd0;\
		conv1_result[0][4][13] <= 18'd0;\
		conv1_result[0][5][0] <= 18'd0;\
		conv1_result[0][5][1] <= 18'd0;\
		conv1_result[0][5][2] <= 18'd0;\
		conv1_result[0][5][3] <= 18'd0;\
		conv1_result[0][5][4] <= 18'd0;\
		conv1_result[0][5][5] <= 18'd0;\
		conv1_result[0][5][6] <= 18'd0;\
		conv1_result[0][5][7] <= 18'd0;\
		conv1_result[0][5][8] <= 18'd0;\
		conv1_result[0][5][9] <= 18'd0;\
		conv1_result[0][5][10] <= 18'd0;\
		conv1_result[0][5][11] <= 18'd0;\
		conv1_result[0][5][12] <= 18'd0;\
		conv1_result[0][5][13] <= 18'd0;\
		conv1_result[0][6][0] <= 18'd0;\
		conv1_result[0][6][1] <= 18'd0;\
		conv1_result[0][6][2] <= 18'd0;\
		conv1_result[0][6][3] <= 18'd0;\
		conv1_result[0][6][4] <= 18'd0;\
		conv1_result[0][6][5] <= 18'd0;\
		conv1_result[0][6][6] <= 18'd0;\
		conv1_result[0][6][7] <= 18'd0;\
		conv1_result[0][6][8] <= 18'd0;\
		conv1_result[0][6][9] <= 18'd0;\
		conv1_result[0][6][10] <= 18'd0;\
		conv1_result[0][6][11] <= 18'd0;\
		conv1_result[0][6][12] <= 18'd0;\
		conv1_result[0][6][13] <= 18'd0;\
		conv1_result[0][7][0] <= 18'd0;\
		conv1_result[0][7][1] <= 18'd0;\
		conv1_result[0][7][2] <= 18'd0;\
		conv1_result[0][7][3] <= 18'd0;\
		conv1_result[0][7][4] <= 18'd0;\
		conv1_result[0][7][5] <= 18'd0;\
		conv1_result[0][7][6] <= 18'd0;\
		conv1_result[0][7][7] <= 18'd0;\
		conv1_result[0][7][8] <= 18'd0;\
		conv1_result[0][7][9] <= 18'd0;\
		conv1_result[0][7][10] <= 18'd0;\
		conv1_result[0][7][11] <= 18'd0;\
		conv1_result[0][7][12] <= 18'd0;\
		conv1_result[0][7][13] <= 18'd0;\
		conv1_result[0][8][0] <= 18'd0;\
		conv1_result[0][8][1] <= 18'd0;\
		conv1_result[0][8][2] <= 18'd0;\
		conv1_result[0][8][3] <= 18'd0;\
		conv1_result[0][8][4] <= 18'd0;\
		conv1_result[0][8][5] <= 18'd0;\
		conv1_result[0][8][6] <= 18'd0;\
		conv1_result[0][8][7] <= 18'd0;\
		conv1_result[0][8][8] <= 18'd0;\
		conv1_result[0][8][9] <= 18'd0;\
		conv1_result[0][8][10] <= 18'd0;\
		conv1_result[0][8][11] <= 18'd0;\
		conv1_result[0][8][12] <= 18'd0;\
		conv1_result[0][8][13] <= 18'd0;\
		conv1_result[0][9][0] <= 18'd0;\
		conv1_result[0][9][1] <= 18'd0;\
		conv1_result[0][9][2] <= 18'd0;\
		conv1_result[0][9][3] <= 18'd0;\
		conv1_result[0][9][4] <= 18'd0;\
		conv1_result[0][9][5] <= 18'd0;\
		conv1_result[0][9][6] <= 18'd0;\
		conv1_result[0][9][7] <= 18'd0;\
		conv1_result[0][9][8] <= 18'd0;\
		conv1_result[0][9][9] <= 18'd0;\
		conv1_result[0][9][10] <= 18'd0;\
		conv1_result[0][9][11] <= 18'd0;\
		conv1_result[0][9][12] <= 18'd0;\
		conv1_result[0][9][13] <= 18'd0;\
		conv1_result[0][10][0] <= 18'd0;\
		conv1_result[0][10][1] <= 18'd0;\
		conv1_result[0][10][2] <= 18'd0;\
		conv1_result[0][10][3] <= 18'd0;\
		conv1_result[0][10][4] <= 18'd0;\
		conv1_result[0][10][5] <= 18'd0;\
		conv1_result[0][10][6] <= 18'd0;\
		conv1_result[0][10][7] <= 18'd0;\
		conv1_result[0][10][8] <= 18'd0;\
		conv1_result[0][10][9] <= 18'd0;\
		conv1_result[0][10][10] <= 18'd0;\
		conv1_result[0][10][11] <= 18'd0;\
		conv1_result[0][10][12] <= 18'd0;\
		conv1_result[0][10][13] <= 18'd0;\
		conv1_result[0][11][0] <= 18'd0;\
		conv1_result[0][11][1] <= 18'd0;\
		conv1_result[0][11][2] <= 18'd0;\
		conv1_result[0][11][3] <= 18'd0;\
		conv1_result[0][11][4] <= 18'd0;\
		conv1_result[0][11][5] <= 18'd0;\
		conv1_result[0][11][6] <= 18'd0;\
		conv1_result[0][11][7] <= 18'd0;\
		conv1_result[0][11][8] <= 18'd0;\
		conv1_result[0][11][9] <= 18'd0;\
		conv1_result[0][11][10] <= 18'd0;\
		conv1_result[0][11][11] <= 18'd0;\
		conv1_result[0][11][12] <= 18'd0;\
		conv1_result[0][11][13] <= 18'd0;\
		conv1_result[0][12][0] <= 18'd0;\
		conv1_result[0][12][1] <= 18'd0;\
		conv1_result[0][12][2] <= 18'd0;\
		conv1_result[0][12][3] <= 18'd0;\
		conv1_result[0][12][4] <= 18'd0;\
		conv1_result[0][12][5] <= 18'd0;\
		conv1_result[0][12][6] <= 18'd0;\
		conv1_result[0][12][7] <= 18'd0;\
		conv1_result[0][12][8] <= 18'd0;\
		conv1_result[0][12][9] <= 18'd0;\
		conv1_result[0][12][10] <= 18'd0;\
		conv1_result[0][12][11] <= 18'd0;\
		conv1_result[0][12][12] <= 18'd0;\
		conv1_result[0][12][13] <= 18'd0;\
		conv1_result[0][13][0] <= 18'd0;\
		conv1_result[0][13][1] <= 18'd0;\
		conv1_result[0][13][2] <= 18'd0;\
		conv1_result[0][13][3] <= 18'd0;\
		conv1_result[0][13][4] <= 18'd0;\
		conv1_result[0][13][5] <= 18'd0;\
		conv1_result[0][13][6] <= 18'd0;\
		conv1_result[0][13][7] <= 18'd0;\
		conv1_result[0][13][8] <= 18'd0;\
		conv1_result[0][13][9] <= 18'd0;\
		conv1_result[0][13][10] <= 18'd0;\
		conv1_result[0][13][11] <= 18'd0;\
		conv1_result[0][13][12] <= 18'd0;\
		conv1_result[0][13][13] <= 18'd0;\
		conv1_result[1][0][0] <= 18'd0;\
		conv1_result[1][0][1] <= 18'd0;\
		conv1_result[1][0][2] <= 18'd0;\
		conv1_result[1][0][3] <= 18'd0;\
		conv1_result[1][0][4] <= 18'd0;\
		conv1_result[1][0][5] <= 18'd0;\
		conv1_result[1][0][6] <= 18'd0;\
		conv1_result[1][0][7] <= 18'd0;\
		conv1_result[1][0][8] <= 18'd0;\
		conv1_result[1][0][9] <= 18'd0;\
		conv1_result[1][0][10] <= 18'd0;\
		conv1_result[1][0][11] <= 18'd0;\
		conv1_result[1][0][12] <= 18'd0;\
		conv1_result[1][0][13] <= 18'd0;\
		conv1_result[1][1][0] <= 18'd0;\
		conv1_result[1][1][1] <= 18'd0;\
		conv1_result[1][1][2] <= 18'd0;\
		conv1_result[1][1][3] <= 18'd0;\
		conv1_result[1][1][4] <= 18'd0;\
		conv1_result[1][1][5] <= 18'd0;\
		conv1_result[1][1][6] <= 18'd0;\
		conv1_result[1][1][7] <= 18'd0;\
		conv1_result[1][1][8] <= 18'd0;\
		conv1_result[1][1][9] <= 18'd0;\
		conv1_result[1][1][10] <= 18'd0;\
		conv1_result[1][1][11] <= 18'd0;\
		conv1_result[1][1][12] <= 18'd0;\
		conv1_result[1][1][13] <= 18'd0;\
		conv1_result[1][2][0] <= 18'd0;\
		conv1_result[1][2][1] <= 18'd0;\
		conv1_result[1][2][2] <= 18'd0;\
		conv1_result[1][2][3] <= 18'd0;\
		conv1_result[1][2][4] <= 18'd0;\
		conv1_result[1][2][5] <= 18'd0;\
		conv1_result[1][2][6] <= 18'd0;\
		conv1_result[1][2][7] <= 18'd0;\
		conv1_result[1][2][8] <= 18'd0;\
		conv1_result[1][2][9] <= 18'd0;\
		conv1_result[1][2][10] <= 18'd0;\
		conv1_result[1][2][11] <= 18'd0;\
		conv1_result[1][2][12] <= 18'd0;\
		conv1_result[1][2][13] <= 18'd0;\
		conv1_result[1][3][0] <= 18'd0;\
		conv1_result[1][3][1] <= 18'd0;\
		conv1_result[1][3][2] <= 18'd0;\
		conv1_result[1][3][3] <= 18'd0;\
		conv1_result[1][3][4] <= 18'd0;\
		conv1_result[1][3][5] <= 18'd0;\
		conv1_result[1][3][6] <= 18'd0;\
		conv1_result[1][3][7] <= 18'd0;\
		conv1_result[1][3][8] <= 18'd0;\
		conv1_result[1][3][9] <= 18'd0;\
		conv1_result[1][3][10] <= 18'd0;\
		conv1_result[1][3][11] <= 18'd0;\
		conv1_result[1][3][12] <= 18'd0;\
		conv1_result[1][3][13] <= 18'd0;\
		conv1_result[1][4][0] <= 18'd0;\
		conv1_result[1][4][1] <= 18'd0;\
		conv1_result[1][4][2] <= 18'd0;\
		conv1_result[1][4][3] <= 18'd0;\
		conv1_result[1][4][4] <= 18'd0;\
		conv1_result[1][4][5] <= 18'd0;\
		conv1_result[1][4][6] <= 18'd0;\
		conv1_result[1][4][7] <= 18'd0;\
		conv1_result[1][4][8] <= 18'd0;\
		conv1_result[1][4][9] <= 18'd0;\
		conv1_result[1][4][10] <= 18'd0;\
		conv1_result[1][4][11] <= 18'd0;\
		conv1_result[1][4][12] <= 18'd0;\
		conv1_result[1][4][13] <= 18'd0;\
		conv1_result[1][5][0] <= 18'd0;\
		conv1_result[1][5][1] <= 18'd0;\
		conv1_result[1][5][2] <= 18'd0;\
		conv1_result[1][5][3] <= 18'd0;\
		conv1_result[1][5][4] <= 18'd0;\
		conv1_result[1][5][5] <= 18'd0;\
		conv1_result[1][5][6] <= 18'd0;\
		conv1_result[1][5][7] <= 18'd0;\
		conv1_result[1][5][8] <= 18'd0;\
		conv1_result[1][5][9] <= 18'd0;\
		conv1_result[1][5][10] <= 18'd0;\
		conv1_result[1][5][11] <= 18'd0;\
		conv1_result[1][5][12] <= 18'd0;\
		conv1_result[1][5][13] <= 18'd0;\
		conv1_result[1][6][0] <= 18'd0;\
		conv1_result[1][6][1] <= 18'd0;\
		conv1_result[1][6][2] <= 18'd0;\
		conv1_result[1][6][3] <= 18'd0;\
		conv1_result[1][6][4] <= 18'd0;\
		conv1_result[1][6][5] <= 18'd0;\
		conv1_result[1][6][6] <= 18'd0;\
		conv1_result[1][6][7] <= 18'd0;\
		conv1_result[1][6][8] <= 18'd0;\
		conv1_result[1][6][9] <= 18'd0;\
		conv1_result[1][6][10] <= 18'd0;\
		conv1_result[1][6][11] <= 18'd0;\
		conv1_result[1][6][12] <= 18'd0;\
		conv1_result[1][6][13] <= 18'd0;\
		conv1_result[1][7][0] <= 18'd0;\
		conv1_result[1][7][1] <= 18'd0;\
		conv1_result[1][7][2] <= 18'd0;\
		conv1_result[1][7][3] <= 18'd0;\
		conv1_result[1][7][4] <= 18'd0;\
		conv1_result[1][7][5] <= 18'd0;\
		conv1_result[1][7][6] <= 18'd0;\
		conv1_result[1][7][7] <= 18'd0;\
		conv1_result[1][7][8] <= 18'd0;\
		conv1_result[1][7][9] <= 18'd0;\
		conv1_result[1][7][10] <= 18'd0;\
		conv1_result[1][7][11] <= 18'd0;\
		conv1_result[1][7][12] <= 18'd0;\
		conv1_result[1][7][13] <= 18'd0;\
		conv1_result[1][8][0] <= 18'd0;\
		conv1_result[1][8][1] <= 18'd0;\
		conv1_result[1][8][2] <= 18'd0;\
		conv1_result[1][8][3] <= 18'd0;\
		conv1_result[1][8][4] <= 18'd0;\
		conv1_result[1][8][5] <= 18'd0;\
		conv1_result[1][8][6] <= 18'd0;\
		conv1_result[1][8][7] <= 18'd0;\
		conv1_result[1][8][8] <= 18'd0;\
		conv1_result[1][8][9] <= 18'd0;\
		conv1_result[1][8][10] <= 18'd0;\
		conv1_result[1][8][11] <= 18'd0;\
		conv1_result[1][8][12] <= 18'd0;\
		conv1_result[1][8][13] <= 18'd0;\
		conv1_result[1][9][0] <= 18'd0;\
		conv1_result[1][9][1] <= 18'd0;\
		conv1_result[1][9][2] <= 18'd0;\
		conv1_result[1][9][3] <= 18'd0;\
		conv1_result[1][9][4] <= 18'd0;\
		conv1_result[1][9][5] <= 18'd0;\
		conv1_result[1][9][6] <= 18'd0;\
		conv1_result[1][9][7] <= 18'd0;\
		conv1_result[1][9][8] <= 18'd0;\
		conv1_result[1][9][9] <= 18'd0;\
		conv1_result[1][9][10] <= 18'd0;\
		conv1_result[1][9][11] <= 18'd0;\
		conv1_result[1][9][12] <= 18'd0;\
		conv1_result[1][9][13] <= 18'd0;\
		conv1_result[1][10][0] <= 18'd0;\
		conv1_result[1][10][1] <= 18'd0;\
		conv1_result[1][10][2] <= 18'd0;\
		conv1_result[1][10][3] <= 18'd0;\
		conv1_result[1][10][4] <= 18'd0;\
		conv1_result[1][10][5] <= 18'd0;\
		conv1_result[1][10][6] <= 18'd0;\
		conv1_result[1][10][7] <= 18'd0;\
		conv1_result[1][10][8] <= 18'd0;\
		conv1_result[1][10][9] <= 18'd0;\
		conv1_result[1][10][10] <= 18'd0;\
		conv1_result[1][10][11] <= 18'd0;\
		conv1_result[1][10][12] <= 18'd0;\
		conv1_result[1][10][13] <= 18'd0;\
		conv1_result[1][11][0] <= 18'd0;\
		conv1_result[1][11][1] <= 18'd0;\
		conv1_result[1][11][2] <= 18'd0;\
		conv1_result[1][11][3] <= 18'd0;\
		conv1_result[1][11][4] <= 18'd0;\
		conv1_result[1][11][5] <= 18'd0;\
		conv1_result[1][11][6] <= 18'd0;\
		conv1_result[1][11][7] <= 18'd0;\
		conv1_result[1][11][8] <= 18'd0;\
		conv1_result[1][11][9] <= 18'd0;\
		conv1_result[1][11][10] <= 18'd0;\
		conv1_result[1][11][11] <= 18'd0;\
		conv1_result[1][11][12] <= 18'd0;\
		conv1_result[1][11][13] <= 18'd0;\
		conv1_result[1][12][0] <= 18'd0;\
		conv1_result[1][12][1] <= 18'd0;\
		conv1_result[1][12][2] <= 18'd0;\
		conv1_result[1][12][3] <= 18'd0;\
		conv1_result[1][12][4] <= 18'd0;\
		conv1_result[1][12][5] <= 18'd0;\
		conv1_result[1][12][6] <= 18'd0;\
		conv1_result[1][12][7] <= 18'd0;\
		conv1_result[1][12][8] <= 18'd0;\
		conv1_result[1][12][9] <= 18'd0;\
		conv1_result[1][12][10] <= 18'd0;\
		conv1_result[1][12][11] <= 18'd0;\
		conv1_result[1][12][12] <= 18'd0;\
		conv1_result[1][12][13] <= 18'd0;\
		conv1_result[1][13][0] <= 18'd0;\
		conv1_result[1][13][1] <= 18'd0;\
		conv1_result[1][13][2] <= 18'd0;\
		conv1_result[1][13][3] <= 18'd0;\
		conv1_result[1][13][4] <= 18'd0;\
		conv1_result[1][13][5] <= 18'd0;\
		conv1_result[1][13][6] <= 18'd0;\
		conv1_result[1][13][7] <= 18'd0;\
		conv1_result[1][13][8] <= 18'd0;\
		conv1_result[1][13][9] <= 18'd0;\
		conv1_result[1][13][10] <= 18'd0;\
		conv1_result[1][13][11] <= 18'd0;\
		conv1_result[1][13][12] <= 18'd0;\
		conv1_result[1][13][13] <= 18'd0;\
		conv1_result[2][0][0] <= 18'd0;\
		conv1_result[2][0][1] <= 18'd0;\
		conv1_result[2][0][2] <= 18'd0;\
		conv1_result[2][0][3] <= 18'd0;\
		conv1_result[2][0][4] <= 18'd0;\
		conv1_result[2][0][5] <= 18'd0;\
		conv1_result[2][0][6] <= 18'd0;\
		conv1_result[2][0][7] <= 18'd0;\
		conv1_result[2][0][8] <= 18'd0;\
		conv1_result[2][0][9] <= 18'd0;\
		conv1_result[2][0][10] <= 18'd0;\
		conv1_result[2][0][11] <= 18'd0;\
		conv1_result[2][0][12] <= 18'd0;\
		conv1_result[2][0][13] <= 18'd0;\
		conv1_result[2][1][0] <= 18'd0;\
		conv1_result[2][1][1] <= 18'd0;\
		conv1_result[2][1][2] <= 18'd0;\
		conv1_result[2][1][3] <= 18'd0;\
		conv1_result[2][1][4] <= 18'd0;\
		conv1_result[2][1][5] <= 18'd0;\
		conv1_result[2][1][6] <= 18'd0;\
		conv1_result[2][1][7] <= 18'd0;\
		conv1_result[2][1][8] <= 18'd0;\
		conv1_result[2][1][9] <= 18'd0;\
		conv1_result[2][1][10] <= 18'd0;\
		conv1_result[2][1][11] <= 18'd0;\
		conv1_result[2][1][12] <= 18'd0;\
		conv1_result[2][1][13] <= 18'd0;\
		conv1_result[2][2][0] <= 18'd0;\
		conv1_result[2][2][1] <= 18'd0;\
		conv1_result[2][2][2] <= 18'd0;\
		conv1_result[2][2][3] <= 18'd0;\
		conv1_result[2][2][4] <= 18'd0;\
		conv1_result[2][2][5] <= 18'd0;\
		conv1_result[2][2][6] <= 18'd0;\
		conv1_result[2][2][7] <= 18'd0;\
		conv1_result[2][2][8] <= 18'd0;\
		conv1_result[2][2][9] <= 18'd0;\
		conv1_result[2][2][10] <= 18'd0;\
		conv1_result[2][2][11] <= 18'd0;\
		conv1_result[2][2][12] <= 18'd0;\
		conv1_result[2][2][13] <= 18'd0;\
		conv1_result[2][3][0] <= 18'd0;\
		conv1_result[2][3][1] <= 18'd0;\
		conv1_result[2][3][2] <= 18'd0;\
		conv1_result[2][3][3] <= 18'd0;\
		conv1_result[2][3][4] <= 18'd0;\
		conv1_result[2][3][5] <= 18'd0;\
		conv1_result[2][3][6] <= 18'd0;\
		conv1_result[2][3][7] <= 18'd0;\
		conv1_result[2][3][8] <= 18'd0;\
		conv1_result[2][3][9] <= 18'd0;\
		conv1_result[2][3][10] <= 18'd0;\
		conv1_result[2][3][11] <= 18'd0;\
		conv1_result[2][3][12] <= 18'd0;\
		conv1_result[2][3][13] <= 18'd0;\
		conv1_result[2][4][0] <= 18'd0;\
		conv1_result[2][4][1] <= 18'd0;\
		conv1_result[2][4][2] <= 18'd0;\
		conv1_result[2][4][3] <= 18'd0;\
		conv1_result[2][4][4] <= 18'd0;\
		conv1_result[2][4][5] <= 18'd0;\
		conv1_result[2][4][6] <= 18'd0;\
		conv1_result[2][4][7] <= 18'd0;\
		conv1_result[2][4][8] <= 18'd0;\
		conv1_result[2][4][9] <= 18'd0;\
		conv1_result[2][4][10] <= 18'd0;\
		conv1_result[2][4][11] <= 18'd0;\
		conv1_result[2][4][12] <= 18'd0;\
		conv1_result[2][4][13] <= 18'd0;\
		conv1_result[2][5][0] <= 18'd0;\
		conv1_result[2][5][1] <= 18'd0;\
		conv1_result[2][5][2] <= 18'd0;\
		conv1_result[2][5][3] <= 18'd0;\
		conv1_result[2][5][4] <= 18'd0;\
		conv1_result[2][5][5] <= 18'd0;\
		conv1_result[2][5][6] <= 18'd0;\
		conv1_result[2][5][7] <= 18'd0;\
		conv1_result[2][5][8] <= 18'd0;\
		conv1_result[2][5][9] <= 18'd0;\
		conv1_result[2][5][10] <= 18'd0;\
		conv1_result[2][5][11] <= 18'd0;\
		conv1_result[2][5][12] <= 18'd0;\
		conv1_result[2][5][13] <= 18'd0;\
		conv1_result[2][6][0] <= 18'd0;\
		conv1_result[2][6][1] <= 18'd0;\
		conv1_result[2][6][2] <= 18'd0;\
		conv1_result[2][6][3] <= 18'd0;\
		conv1_result[2][6][4] <= 18'd0;\
		conv1_result[2][6][5] <= 18'd0;\
		conv1_result[2][6][6] <= 18'd0;\
		conv1_result[2][6][7] <= 18'd0;\
		conv1_result[2][6][8] <= 18'd0;\
		conv1_result[2][6][9] <= 18'd0;\
		conv1_result[2][6][10] <= 18'd0;\
		conv1_result[2][6][11] <= 18'd0;\
		conv1_result[2][6][12] <= 18'd0;\
		conv1_result[2][6][13] <= 18'd0;\
		conv1_result[2][7][0] <= 18'd0;\
		conv1_result[2][7][1] <= 18'd0;\
		conv1_result[2][7][2] <= 18'd0;\
		conv1_result[2][7][3] <= 18'd0;\
		conv1_result[2][7][4] <= 18'd0;\
		conv1_result[2][7][5] <= 18'd0;\
		conv1_result[2][7][6] <= 18'd0;\
		conv1_result[2][7][7] <= 18'd0;\
		conv1_result[2][7][8] <= 18'd0;\
		conv1_result[2][7][9] <= 18'd0;\
		conv1_result[2][7][10] <= 18'd0;\
		conv1_result[2][7][11] <= 18'd0;\
		conv1_result[2][7][12] <= 18'd0;\
		conv1_result[2][7][13] <= 18'd0;\
		conv1_result[2][8][0] <= 18'd0;\
		conv1_result[2][8][1] <= 18'd0;\
		conv1_result[2][8][2] <= 18'd0;\
		conv1_result[2][8][3] <= 18'd0;\
		conv1_result[2][8][4] <= 18'd0;\
		conv1_result[2][8][5] <= 18'd0;\
		conv1_result[2][8][6] <= 18'd0;\
		conv1_result[2][8][7] <= 18'd0;\
		conv1_result[2][8][8] <= 18'd0;\
		conv1_result[2][8][9] <= 18'd0;\
		conv1_result[2][8][10] <= 18'd0;\
		conv1_result[2][8][11] <= 18'd0;\
		conv1_result[2][8][12] <= 18'd0;\
		conv1_result[2][8][13] <= 18'd0;\
		conv1_result[2][9][0] <= 18'd0;\
		conv1_result[2][9][1] <= 18'd0;\
		conv1_result[2][9][2] <= 18'd0;\
		conv1_result[2][9][3] <= 18'd0;\
		conv1_result[2][9][4] <= 18'd0;\
		conv1_result[2][9][5] <= 18'd0;\
		conv1_result[2][9][6] <= 18'd0;\
		conv1_result[2][9][7] <= 18'd0;\
		conv1_result[2][9][8] <= 18'd0;\
		conv1_result[2][9][9] <= 18'd0;\
		conv1_result[2][9][10] <= 18'd0;\
		conv1_result[2][9][11] <= 18'd0;\
		conv1_result[2][9][12] <= 18'd0;\
		conv1_result[2][9][13] <= 18'd0;\
		conv1_result[2][10][0] <= 18'd0;\
		conv1_result[2][10][1] <= 18'd0;\
		conv1_result[2][10][2] <= 18'd0;\
		conv1_result[2][10][3] <= 18'd0;\
		conv1_result[2][10][4] <= 18'd0;\
		conv1_result[2][10][5] <= 18'd0;\
		conv1_result[2][10][6] <= 18'd0;\
		conv1_result[2][10][7] <= 18'd0;\
		conv1_result[2][10][8] <= 18'd0;\
		conv1_result[2][10][9] <= 18'd0;\
		conv1_result[2][10][10] <= 18'd0;\
		conv1_result[2][10][11] <= 18'd0;\
		conv1_result[2][10][12] <= 18'd0;\
		conv1_result[2][10][13] <= 18'd0;\
		conv1_result[2][11][0] <= 18'd0;\
		conv1_result[2][11][1] <= 18'd0;\
		conv1_result[2][11][2] <= 18'd0;\
		conv1_result[2][11][3] <= 18'd0;\
		conv1_result[2][11][4] <= 18'd0;\
		conv1_result[2][11][5] <= 18'd0;\
		conv1_result[2][11][6] <= 18'd0;\
		conv1_result[2][11][7] <= 18'd0;\
		conv1_result[2][11][8] <= 18'd0;\
		conv1_result[2][11][9] <= 18'd0;\
		conv1_result[2][11][10] <= 18'd0;\
		conv1_result[2][11][11] <= 18'd0;\
		conv1_result[2][11][12] <= 18'd0;\
		conv1_result[2][11][13] <= 18'd0;\
		conv1_result[2][12][0] <= 18'd0;\
		conv1_result[2][12][1] <= 18'd0;\
		conv1_result[2][12][2] <= 18'd0;\
		conv1_result[2][12][3] <= 18'd0;\
		conv1_result[2][12][4] <= 18'd0;\
		conv1_result[2][12][5] <= 18'd0;\
		conv1_result[2][12][6] <= 18'd0;\
		conv1_result[2][12][7] <= 18'd0;\
		conv1_result[2][12][8] <= 18'd0;\
		conv1_result[2][12][9] <= 18'd0;\
		conv1_result[2][12][10] <= 18'd0;\
		conv1_result[2][12][11] <= 18'd0;\
		conv1_result[2][12][12] <= 18'd0;\
		conv1_result[2][12][13] <= 18'd0;\
		conv1_result[2][13][0] <= 18'd0;\
		conv1_result[2][13][1] <= 18'd0;\
		conv1_result[2][13][2] <= 18'd0;\
		conv1_result[2][13][3] <= 18'd0;\
		conv1_result[2][13][4] <= 18'd0;\
		conv1_result[2][13][5] <= 18'd0;\
		conv1_result[2][13][6] <= 18'd0;\
		conv1_result[2][13][7] <= 18'd0;\
		conv1_result[2][13][8] <= 18'd0;\
		conv1_result[2][13][9] <= 18'd0;\
		conv1_result[2][13][10] <= 18'd0;\
		conv1_result[2][13][11] <= 18'd0;\
		conv1_result[2][13][12] <= 18'd0;\
		conv1_result[2][13][13] <= 18'd0;\
		conv1_result[3][0][0] <= 18'd0;\
		conv1_result[3][0][1] <= 18'd0;\
		conv1_result[3][0][2] <= 18'd0;\
		conv1_result[3][0][3] <= 18'd0;\
		conv1_result[3][0][4] <= 18'd0;\
		conv1_result[3][0][5] <= 18'd0;\
		conv1_result[3][0][6] <= 18'd0;\
		conv1_result[3][0][7] <= 18'd0;\
		conv1_result[3][0][8] <= 18'd0;\
		conv1_result[3][0][9] <= 18'd0;\
		conv1_result[3][0][10] <= 18'd0;\
		conv1_result[3][0][11] <= 18'd0;\
		conv1_result[3][0][12] <= 18'd0;\
		conv1_result[3][0][13] <= 18'd0;\
		conv1_result[3][1][0] <= 18'd0;\
		conv1_result[3][1][1] <= 18'd0;\
		conv1_result[3][1][2] <= 18'd0;\
		conv1_result[3][1][3] <= 18'd0;\
		conv1_result[3][1][4] <= 18'd0;\
		conv1_result[3][1][5] <= 18'd0;\
		conv1_result[3][1][6] <= 18'd0;\
		conv1_result[3][1][7] <= 18'd0;\
		conv1_result[3][1][8] <= 18'd0;\
		conv1_result[3][1][9] <= 18'd0;\
		conv1_result[3][1][10] <= 18'd0;\
		conv1_result[3][1][11] <= 18'd0;\
		conv1_result[3][1][12] <= 18'd0;\
		conv1_result[3][1][13] <= 18'd0;\
		conv1_result[3][2][0] <= 18'd0;\
		conv1_result[3][2][1] <= 18'd0;\
		conv1_result[3][2][2] <= 18'd0;\
		conv1_result[3][2][3] <= 18'd0;\
		conv1_result[3][2][4] <= 18'd0;\
		conv1_result[3][2][5] <= 18'd0;\
		conv1_result[3][2][6] <= 18'd0;\
		conv1_result[3][2][7] <= 18'd0;\
		conv1_result[3][2][8] <= 18'd0;\
		conv1_result[3][2][9] <= 18'd0;\
		conv1_result[3][2][10] <= 18'd0;\
		conv1_result[3][2][11] <= 18'd0;\
		conv1_result[3][2][12] <= 18'd0;\
		conv1_result[3][2][13] <= 18'd0;\
		conv1_result[3][3][0] <= 18'd0;\
		conv1_result[3][3][1] <= 18'd0;\
		conv1_result[3][3][2] <= 18'd0;\
		conv1_result[3][3][3] <= 18'd0;\
		conv1_result[3][3][4] <= 18'd0;\
		conv1_result[3][3][5] <= 18'd0;\
		conv1_result[3][3][6] <= 18'd0;\
		conv1_result[3][3][7] <= 18'd0;\
		conv1_result[3][3][8] <= 18'd0;\
		conv1_result[3][3][9] <= 18'd0;\
		conv1_result[3][3][10] <= 18'd0;\
		conv1_result[3][3][11] <= 18'd0;\
		conv1_result[3][3][12] <= 18'd0;\
		conv1_result[3][3][13] <= 18'd0;\
		conv1_result[3][4][0] <= 18'd0;\
		conv1_result[3][4][1] <= 18'd0;\
		conv1_result[3][4][2] <= 18'd0;\
		conv1_result[3][4][3] <= 18'd0;\
		conv1_result[3][4][4] <= 18'd0;\
		conv1_result[3][4][5] <= 18'd0;\
		conv1_result[3][4][6] <= 18'd0;\
		conv1_result[3][4][7] <= 18'd0;\
		conv1_result[3][4][8] <= 18'd0;\
		conv1_result[3][4][9] <= 18'd0;\
		conv1_result[3][4][10] <= 18'd0;\
		conv1_result[3][4][11] <= 18'd0;\
		conv1_result[3][4][12] <= 18'd0;\
		conv1_result[3][4][13] <= 18'd0;\
		conv1_result[3][5][0] <= 18'd0;\
		conv1_result[3][5][1] <= 18'd0;\
		conv1_result[3][5][2] <= 18'd0;\
		conv1_result[3][5][3] <= 18'd0;\
		conv1_result[3][5][4] <= 18'd0;\
		conv1_result[3][5][5] <= 18'd0;\
		conv1_result[3][5][6] <= 18'd0;\
		conv1_result[3][5][7] <= 18'd0;\
		conv1_result[3][5][8] <= 18'd0;\
		conv1_result[3][5][9] <= 18'd0;\
		conv1_result[3][5][10] <= 18'd0;\
		conv1_result[3][5][11] <= 18'd0;\
		conv1_result[3][5][12] <= 18'd0;\
		conv1_result[3][5][13] <= 18'd0;\
		conv1_result[3][6][0] <= 18'd0;\
		conv1_result[3][6][1] <= 18'd0;\
		conv1_result[3][6][2] <= 18'd0;\
		conv1_result[3][6][3] <= 18'd0;\
		conv1_result[3][6][4] <= 18'd0;\
		conv1_result[3][6][5] <= 18'd0;\
		conv1_result[3][6][6] <= 18'd0;\
		conv1_result[3][6][7] <= 18'd0;\
		conv1_result[3][6][8] <= 18'd0;\
		conv1_result[3][6][9] <= 18'd0;\
		conv1_result[3][6][10] <= 18'd0;\
		conv1_result[3][6][11] <= 18'd0;\
		conv1_result[3][6][12] <= 18'd0;\
		conv1_result[3][6][13] <= 18'd0;\
		conv1_result[3][7][0] <= 18'd0;\
		conv1_result[3][7][1] <= 18'd0;\
		conv1_result[3][7][2] <= 18'd0;\
		conv1_result[3][7][3] <= 18'd0;\
		conv1_result[3][7][4] <= 18'd0;\
		conv1_result[3][7][5] <= 18'd0;\
		conv1_result[3][7][6] <= 18'd0;\
		conv1_result[3][7][7] <= 18'd0;\
		conv1_result[3][7][8] <= 18'd0;\
		conv1_result[3][7][9] <= 18'd0;\
		conv1_result[3][7][10] <= 18'd0;\
		conv1_result[3][7][11] <= 18'd0;\
		conv1_result[3][7][12] <= 18'd0;\
		conv1_result[3][7][13] <= 18'd0;\
		conv1_result[3][8][0] <= 18'd0;\
		conv1_result[3][8][1] <= 18'd0;\
		conv1_result[3][8][2] <= 18'd0;\
		conv1_result[3][8][3] <= 18'd0;\
		conv1_result[3][8][4] <= 18'd0;\
		conv1_result[3][8][5] <= 18'd0;\
		conv1_result[3][8][6] <= 18'd0;\
		conv1_result[3][8][7] <= 18'd0;\
		conv1_result[3][8][8] <= 18'd0;\
		conv1_result[3][8][9] <= 18'd0;\
		conv1_result[3][8][10] <= 18'd0;\
		conv1_result[3][8][11] <= 18'd0;\
		conv1_result[3][8][12] <= 18'd0;\
		conv1_result[3][8][13] <= 18'd0;\
		conv1_result[3][9][0] <= 18'd0;\
		conv1_result[3][9][1] <= 18'd0;\
		conv1_result[3][9][2] <= 18'd0;\
		conv1_result[3][9][3] <= 18'd0;\
		conv1_result[3][9][4] <= 18'd0;\
		conv1_result[3][9][5] <= 18'd0;\
		conv1_result[3][9][6] <= 18'd0;\
		conv1_result[3][9][7] <= 18'd0;\
		conv1_result[3][9][8] <= 18'd0;\
		conv1_result[3][9][9] <= 18'd0;\
		conv1_result[3][9][10] <= 18'd0;\
		conv1_result[3][9][11] <= 18'd0;\
		conv1_result[3][9][12] <= 18'd0;\
		conv1_result[3][9][13] <= 18'd0;\
		conv1_result[3][10][0] <= 18'd0;\
		conv1_result[3][10][1] <= 18'd0;\
		conv1_result[3][10][2] <= 18'd0;\
		conv1_result[3][10][3] <= 18'd0;\
		conv1_result[3][10][4] <= 18'd0;\
		conv1_result[3][10][5] <= 18'd0;\
		conv1_result[3][10][6] <= 18'd0;\
		conv1_result[3][10][7] <= 18'd0;\
		conv1_result[3][10][8] <= 18'd0;\
		conv1_result[3][10][9] <= 18'd0;\
		conv1_result[3][10][10] <= 18'd0;\
		conv1_result[3][10][11] <= 18'd0;\
		conv1_result[3][10][12] <= 18'd0;\
		conv1_result[3][10][13] <= 18'd0;\
		conv1_result[3][11][0] <= 18'd0;\
		conv1_result[3][11][1] <= 18'd0;\
		conv1_result[3][11][2] <= 18'd0;\
		conv1_result[3][11][3] <= 18'd0;\
		conv1_result[3][11][4] <= 18'd0;\
		conv1_result[3][11][5] <= 18'd0;\
		conv1_result[3][11][6] <= 18'd0;\
		conv1_result[3][11][7] <= 18'd0;\
		conv1_result[3][11][8] <= 18'd0;\
		conv1_result[3][11][9] <= 18'd0;\
		conv1_result[3][11][10] <= 18'd0;\
		conv1_result[3][11][11] <= 18'd0;\
		conv1_result[3][11][12] <= 18'd0;\
		conv1_result[3][11][13] <= 18'd0;\
		conv1_result[3][12][0] <= 18'd0;\
		conv1_result[3][12][1] <= 18'd0;\
		conv1_result[3][12][2] <= 18'd0;\
		conv1_result[3][12][3] <= 18'd0;\
		conv1_result[3][12][4] <= 18'd0;\
		conv1_result[3][12][5] <= 18'd0;\
		conv1_result[3][12][6] <= 18'd0;\
		conv1_result[3][12][7] <= 18'd0;\
		conv1_result[3][12][8] <= 18'd0;\
		conv1_result[3][12][9] <= 18'd0;\
		conv1_result[3][12][10] <= 18'd0;\
		conv1_result[3][12][11] <= 18'd0;\
		conv1_result[3][12][12] <= 18'd0;\
		conv1_result[3][12][13] <= 18'd0;\
		conv1_result[3][13][0] <= 18'd0;\
		conv1_result[3][13][1] <= 18'd0;\
		conv1_result[3][13][2] <= 18'd0;\
		conv1_result[3][13][3] <= 18'd0;\
		conv1_result[3][13][4] <= 18'd0;\
		conv1_result[3][13][5] <= 18'd0;\
		conv1_result[3][13][6] <= 18'd0;\
		conv1_result[3][13][7] <= 18'd0;\
		conv1_result[3][13][8] <= 18'd0;\
		conv1_result[3][13][9] <= 18'd0;\
		conv1_result[3][13][10] <= 18'd0;\
		conv1_result[3][13][11] <= 18'd0;\
		conv1_result[3][13][12] <= 18'd0;\
		conv1_result[3][13][13] <= 18'd0;\
		conv1_result[4][0][0] <= 18'd0;\
		conv1_result[4][0][1] <= 18'd0;\
		conv1_result[4][0][2] <= 18'd0;\
		conv1_result[4][0][3] <= 18'd0;\
		conv1_result[4][0][4] <= 18'd0;\
		conv1_result[4][0][5] <= 18'd0;\
		conv1_result[4][0][6] <= 18'd0;\
		conv1_result[4][0][7] <= 18'd0;\
		conv1_result[4][0][8] <= 18'd0;\
		conv1_result[4][0][9] <= 18'd0;\
		conv1_result[4][0][10] <= 18'd0;\
		conv1_result[4][0][11] <= 18'd0;\
		conv1_result[4][0][12] <= 18'd0;\
		conv1_result[4][0][13] <= 18'd0;\
		conv1_result[4][1][0] <= 18'd0;\
		conv1_result[4][1][1] <= 18'd0;\
		conv1_result[4][1][2] <= 18'd0;\
		conv1_result[4][1][3] <= 18'd0;\
		conv1_result[4][1][4] <= 18'd0;\
		conv1_result[4][1][5] <= 18'd0;\
		conv1_result[4][1][6] <= 18'd0;\
		conv1_result[4][1][7] <= 18'd0;\
		conv1_result[4][1][8] <= 18'd0;\
		conv1_result[4][1][9] <= 18'd0;\
		conv1_result[4][1][10] <= 18'd0;\
		conv1_result[4][1][11] <= 18'd0;\
		conv1_result[4][1][12] <= 18'd0;\
		conv1_result[4][1][13] <= 18'd0;\
		conv1_result[4][2][0] <= 18'd0;\
		conv1_result[4][2][1] <= 18'd0;\
		conv1_result[4][2][2] <= 18'd0;\
		conv1_result[4][2][3] <= 18'd0;\
		conv1_result[4][2][4] <= 18'd0;\
		conv1_result[4][2][5] <= 18'd0;\
		conv1_result[4][2][6] <= 18'd0;\
		conv1_result[4][2][7] <= 18'd0;\
		conv1_result[4][2][8] <= 18'd0;\
		conv1_result[4][2][9] <= 18'd0;\
		conv1_result[4][2][10] <= 18'd0;\
		conv1_result[4][2][11] <= 18'd0;\
		conv1_result[4][2][12] <= 18'd0;\
		conv1_result[4][2][13] <= 18'd0;\
		conv1_result[4][3][0] <= 18'd0;\
		conv1_result[4][3][1] <= 18'd0;\
		conv1_result[4][3][2] <= 18'd0;\
		conv1_result[4][3][3] <= 18'd0;\
		conv1_result[4][3][4] <= 18'd0;\
		conv1_result[4][3][5] <= 18'd0;\
		conv1_result[4][3][6] <= 18'd0;\
		conv1_result[4][3][7] <= 18'd0;\
		conv1_result[4][3][8] <= 18'd0;\
		conv1_result[4][3][9] <= 18'd0;\
		conv1_result[4][3][10] <= 18'd0;\
		conv1_result[4][3][11] <= 18'd0;\
		conv1_result[4][3][12] <= 18'd0;\
		conv1_result[4][3][13] <= 18'd0;\
		conv1_result[4][4][0] <= 18'd0;\
		conv1_result[4][4][1] <= 18'd0;\
		conv1_result[4][4][2] <= 18'd0;\
		conv1_result[4][4][3] <= 18'd0;\
		conv1_result[4][4][4] <= 18'd0;\
		conv1_result[4][4][5] <= 18'd0;\
		conv1_result[4][4][6] <= 18'd0;\
		conv1_result[4][4][7] <= 18'd0;\
		conv1_result[4][4][8] <= 18'd0;\
		conv1_result[4][4][9] <= 18'd0;\
		conv1_result[4][4][10] <= 18'd0;\
		conv1_result[4][4][11] <= 18'd0;\
		conv1_result[4][4][12] <= 18'd0;\
		conv1_result[4][4][13] <= 18'd0;\
		conv1_result[4][5][0] <= 18'd0;\
		conv1_result[4][5][1] <= 18'd0;\
		conv1_result[4][5][2] <= 18'd0;\
		conv1_result[4][5][3] <= 18'd0;\
		conv1_result[4][5][4] <= 18'd0;\
		conv1_result[4][5][5] <= 18'd0;\
		conv1_result[4][5][6] <= 18'd0;\
		conv1_result[4][5][7] <= 18'd0;\
		conv1_result[4][5][8] <= 18'd0;\
		conv1_result[4][5][9] <= 18'd0;\
		conv1_result[4][5][10] <= 18'd0;\
		conv1_result[4][5][11] <= 18'd0;\
		conv1_result[4][5][12] <= 18'd0;\
		conv1_result[4][5][13] <= 18'd0;\
		conv1_result[4][6][0] <= 18'd0;\
		conv1_result[4][6][1] <= 18'd0;\
		conv1_result[4][6][2] <= 18'd0;\
		conv1_result[4][6][3] <= 18'd0;\
		conv1_result[4][6][4] <= 18'd0;\
		conv1_result[4][6][5] <= 18'd0;\
		conv1_result[4][6][6] <= 18'd0;\
		conv1_result[4][6][7] <= 18'd0;\
		conv1_result[4][6][8] <= 18'd0;\
		conv1_result[4][6][9] <= 18'd0;\
		conv1_result[4][6][10] <= 18'd0;\
		conv1_result[4][6][11] <= 18'd0;\
		conv1_result[4][6][12] <= 18'd0;\
		conv1_result[4][6][13] <= 18'd0;\
		conv1_result[4][7][0] <= 18'd0;\
		conv1_result[4][7][1] <= 18'd0;\
		conv1_result[4][7][2] <= 18'd0;\
		conv1_result[4][7][3] <= 18'd0;\
		conv1_result[4][7][4] <= 18'd0;\
		conv1_result[4][7][5] <= 18'd0;\
		conv1_result[4][7][6] <= 18'd0;\
		conv1_result[4][7][7] <= 18'd0;\
		conv1_result[4][7][8] <= 18'd0;\
		conv1_result[4][7][9] <= 18'd0;\
		conv1_result[4][7][10] <= 18'd0;\
		conv1_result[4][7][11] <= 18'd0;\
		conv1_result[4][7][12] <= 18'd0;\
		conv1_result[4][7][13] <= 18'd0;\
		conv1_result[4][8][0] <= 18'd0;\
		conv1_result[4][8][1] <= 18'd0;\
		conv1_result[4][8][2] <= 18'd0;\
		conv1_result[4][8][3] <= 18'd0;\
		conv1_result[4][8][4] <= 18'd0;\
		conv1_result[4][8][5] <= 18'd0;\
		conv1_result[4][8][6] <= 18'd0;\
		conv1_result[4][8][7] <= 18'd0;\
		conv1_result[4][8][8] <= 18'd0;\
		conv1_result[4][8][9] <= 18'd0;\
		conv1_result[4][8][10] <= 18'd0;\
		conv1_result[4][8][11] <= 18'd0;\
		conv1_result[4][8][12] <= 18'd0;\
		conv1_result[4][8][13] <= 18'd0;\
		conv1_result[4][9][0] <= 18'd0;\
		conv1_result[4][9][1] <= 18'd0;\
		conv1_result[4][9][2] <= 18'd0;\
		conv1_result[4][9][3] <= 18'd0;\
		conv1_result[4][9][4] <= 18'd0;\
		conv1_result[4][9][5] <= 18'd0;\
		conv1_result[4][9][6] <= 18'd0;\
		conv1_result[4][9][7] <= 18'd0;\
		conv1_result[4][9][8] <= 18'd0;\
		conv1_result[4][9][9] <= 18'd0;\
		conv1_result[4][9][10] <= 18'd0;\
		conv1_result[4][9][11] <= 18'd0;\
		conv1_result[4][9][12] <= 18'd0;\
		conv1_result[4][9][13] <= 18'd0;\
		conv1_result[4][10][0] <= 18'd0;\
		conv1_result[4][10][1] <= 18'd0;\
		conv1_result[4][10][2] <= 18'd0;\
		conv1_result[4][10][3] <= 18'd0;\
		conv1_result[4][10][4] <= 18'd0;\
		conv1_result[4][10][5] <= 18'd0;\
		conv1_result[4][10][6] <= 18'd0;\
		conv1_result[4][10][7] <= 18'd0;\
		conv1_result[4][10][8] <= 18'd0;\
		conv1_result[4][10][9] <= 18'd0;\
		conv1_result[4][10][10] <= 18'd0;\
		conv1_result[4][10][11] <= 18'd0;\
		conv1_result[4][10][12] <= 18'd0;\
		conv1_result[4][10][13] <= 18'd0;\
		conv1_result[4][11][0] <= 18'd0;\
		conv1_result[4][11][1] <= 18'd0;\
		conv1_result[4][11][2] <= 18'd0;\
		conv1_result[4][11][3] <= 18'd0;\
		conv1_result[4][11][4] <= 18'd0;\
		conv1_result[4][11][5] <= 18'd0;\
		conv1_result[4][11][6] <= 18'd0;\
		conv1_result[4][11][7] <= 18'd0;\
		conv1_result[4][11][8] <= 18'd0;\
		conv1_result[4][11][9] <= 18'd0;\
		conv1_result[4][11][10] <= 18'd0;\
		conv1_result[4][11][11] <= 18'd0;\
		conv1_result[4][11][12] <= 18'd0;\
		conv1_result[4][11][13] <= 18'd0;\
		conv1_result[4][12][0] <= 18'd0;\
		conv1_result[4][12][1] <= 18'd0;\
		conv1_result[4][12][2] <= 18'd0;\
		conv1_result[4][12][3] <= 18'd0;\
		conv1_result[4][12][4] <= 18'd0;\
		conv1_result[4][12][5] <= 18'd0;\
		conv1_result[4][12][6] <= 18'd0;\
		conv1_result[4][12][7] <= 18'd0;\
		conv1_result[4][12][8] <= 18'd0;\
		conv1_result[4][12][9] <= 18'd0;\
		conv1_result[4][12][10] <= 18'd0;\
		conv1_result[4][12][11] <= 18'd0;\
		conv1_result[4][12][12] <= 18'd0;\
		conv1_result[4][12][13] <= 18'd0;\
		conv1_result[4][13][0] <= 18'd0;\
		conv1_result[4][13][1] <= 18'd0;\
		conv1_result[4][13][2] <= 18'd0;\
		conv1_result[4][13][3] <= 18'd0;\
		conv1_result[4][13][4] <= 18'd0;\
		conv1_result[4][13][5] <= 18'd0;\
		conv1_result[4][13][6] <= 18'd0;\
		conv1_result[4][13][7] <= 18'd0;\
		conv1_result[4][13][8] <= 18'd0;\
		conv1_result[4][13][9] <= 18'd0;\
		conv1_result[4][13][10] <= 18'd0;\
		conv1_result[4][13][11] <= 18'd0;\
		conv1_result[4][13][12] <= 18'd0;\
		conv1_result[4][13][13] <= 18'd0;\
		conv1_result[5][0][0] <= 18'd0;\
		conv1_result[5][0][1] <= 18'd0;\
		conv1_result[5][0][2] <= 18'd0;\
		conv1_result[5][0][3] <= 18'd0;\
		conv1_result[5][0][4] <= 18'd0;\
		conv1_result[5][0][5] <= 18'd0;\
		conv1_result[5][0][6] <= 18'd0;\
		conv1_result[5][0][7] <= 18'd0;\
		conv1_result[5][0][8] <= 18'd0;\
		conv1_result[5][0][9] <= 18'd0;\
		conv1_result[5][0][10] <= 18'd0;\
		conv1_result[5][0][11] <= 18'd0;\
		conv1_result[5][0][12] <= 18'd0;\
		conv1_result[5][0][13] <= 18'd0;\
		conv1_result[5][1][0] <= 18'd0;\
		conv1_result[5][1][1] <= 18'd0;\
		conv1_result[5][1][2] <= 18'd0;\
		conv1_result[5][1][3] <= 18'd0;\
		conv1_result[5][1][4] <= 18'd0;\
		conv1_result[5][1][5] <= 18'd0;\
		conv1_result[5][1][6] <= 18'd0;\
		conv1_result[5][1][7] <= 18'd0;\
		conv1_result[5][1][8] <= 18'd0;\
		conv1_result[5][1][9] <= 18'd0;\
		conv1_result[5][1][10] <= 18'd0;\
		conv1_result[5][1][11] <= 18'd0;\
		conv1_result[5][1][12] <= 18'd0;\
		conv1_result[5][1][13] <= 18'd0;\
		conv1_result[5][2][0] <= 18'd0;\
		conv1_result[5][2][1] <= 18'd0;\
		conv1_result[5][2][2] <= 18'd0;\
		conv1_result[5][2][3] <= 18'd0;\
		conv1_result[5][2][4] <= 18'd0;\
		conv1_result[5][2][5] <= 18'd0;\
		conv1_result[5][2][6] <= 18'd0;\
		conv1_result[5][2][7] <= 18'd0;\
		conv1_result[5][2][8] <= 18'd0;\
		conv1_result[5][2][9] <= 18'd0;\
		conv1_result[5][2][10] <= 18'd0;\
		conv1_result[5][2][11] <= 18'd0;\
		conv1_result[5][2][12] <= 18'd0;\
		conv1_result[5][2][13] <= 18'd0;\
		conv1_result[5][3][0] <= 18'd0;\
		conv1_result[5][3][1] <= 18'd0;\
		conv1_result[5][3][2] <= 18'd0;\
		conv1_result[5][3][3] <= 18'd0;\
		conv1_result[5][3][4] <= 18'd0;\
		conv1_result[5][3][5] <= 18'd0;\
		conv1_result[5][3][6] <= 18'd0;\
		conv1_result[5][3][7] <= 18'd0;\
		conv1_result[5][3][8] <= 18'd0;\
		conv1_result[5][3][9] <= 18'd0;\
		conv1_result[5][3][10] <= 18'd0;\
		conv1_result[5][3][11] <= 18'd0;\
		conv1_result[5][3][12] <= 18'd0;\
		conv1_result[5][3][13] <= 18'd0;\
		conv1_result[5][4][0] <= 18'd0;\
		conv1_result[5][4][1] <= 18'd0;\
		conv1_result[5][4][2] <= 18'd0;\
		conv1_result[5][4][3] <= 18'd0;\
		conv1_result[5][4][4] <= 18'd0;\
		conv1_result[5][4][5] <= 18'd0;\
		conv1_result[5][4][6] <= 18'd0;\
		conv1_result[5][4][7] <= 18'd0;\
		conv1_result[5][4][8] <= 18'd0;\
		conv1_result[5][4][9] <= 18'd0;\
		conv1_result[5][4][10] <= 18'd0;\
		conv1_result[5][4][11] <= 18'd0;\
		conv1_result[5][4][12] <= 18'd0;\
		conv1_result[5][4][13] <= 18'd0;\
		conv1_result[5][5][0] <= 18'd0;\
		conv1_result[5][5][1] <= 18'd0;\
		conv1_result[5][5][2] <= 18'd0;\
		conv1_result[5][5][3] <= 18'd0;\
		conv1_result[5][5][4] <= 18'd0;\
		conv1_result[5][5][5] <= 18'd0;\
		conv1_result[5][5][6] <= 18'd0;\
		conv1_result[5][5][7] <= 18'd0;\
		conv1_result[5][5][8] <= 18'd0;\
		conv1_result[5][5][9] <= 18'd0;\
		conv1_result[5][5][10] <= 18'd0;\
		conv1_result[5][5][11] <= 18'd0;\
		conv1_result[5][5][12] <= 18'd0;\
		conv1_result[5][5][13] <= 18'd0;\
		conv1_result[5][6][0] <= 18'd0;\
		conv1_result[5][6][1] <= 18'd0;\
		conv1_result[5][6][2] <= 18'd0;\
		conv1_result[5][6][3] <= 18'd0;\
		conv1_result[5][6][4] <= 18'd0;\
		conv1_result[5][6][5] <= 18'd0;\
		conv1_result[5][6][6] <= 18'd0;\
		conv1_result[5][6][7] <= 18'd0;\
		conv1_result[5][6][8] <= 18'd0;\
		conv1_result[5][6][9] <= 18'd0;\
		conv1_result[5][6][10] <= 18'd0;\
		conv1_result[5][6][11] <= 18'd0;\
		conv1_result[5][6][12] <= 18'd0;\
		conv1_result[5][6][13] <= 18'd0;\
		conv1_result[5][7][0] <= 18'd0;\
		conv1_result[5][7][1] <= 18'd0;\
		conv1_result[5][7][2] <= 18'd0;\
		conv1_result[5][7][3] <= 18'd0;\
		conv1_result[5][7][4] <= 18'd0;\
		conv1_result[5][7][5] <= 18'd0;\
		conv1_result[5][7][6] <= 18'd0;\
		conv1_result[5][7][7] <= 18'd0;\
		conv1_result[5][7][8] <= 18'd0;\
		conv1_result[5][7][9] <= 18'd0;\
		conv1_result[5][7][10] <= 18'd0;\
		conv1_result[5][7][11] <= 18'd0;\
		conv1_result[5][7][12] <= 18'd0;\
		conv1_result[5][7][13] <= 18'd0;\
		conv1_result[5][8][0] <= 18'd0;\
		conv1_result[5][8][1] <= 18'd0;\
		conv1_result[5][8][2] <= 18'd0;\
		conv1_result[5][8][3] <= 18'd0;\
		conv1_result[5][8][4] <= 18'd0;\
		conv1_result[5][8][5] <= 18'd0;\
		conv1_result[5][8][6] <= 18'd0;\
		conv1_result[5][8][7] <= 18'd0;\
		conv1_result[5][8][8] <= 18'd0;\
		conv1_result[5][8][9] <= 18'd0;\
		conv1_result[5][8][10] <= 18'd0;\
		conv1_result[5][8][11] <= 18'd0;\
		conv1_result[5][8][12] <= 18'd0;\
		conv1_result[5][8][13] <= 18'd0;\
		conv1_result[5][9][0] <= 18'd0;\
		conv1_result[5][9][1] <= 18'd0;\
		conv1_result[5][9][2] <= 18'd0;\
		conv1_result[5][9][3] <= 18'd0;\
		conv1_result[5][9][4] <= 18'd0;\
		conv1_result[5][9][5] <= 18'd0;\
		conv1_result[5][9][6] <= 18'd0;\
		conv1_result[5][9][7] <= 18'd0;\
		conv1_result[5][9][8] <= 18'd0;\
		conv1_result[5][9][9] <= 18'd0;\
		conv1_result[5][9][10] <= 18'd0;\
		conv1_result[5][9][11] <= 18'd0;\
		conv1_result[5][9][12] <= 18'd0;\
		conv1_result[5][9][13] <= 18'd0;\
		conv1_result[5][10][0] <= 18'd0;\
		conv1_result[5][10][1] <= 18'd0;\
		conv1_result[5][10][2] <= 18'd0;\
		conv1_result[5][10][3] <= 18'd0;\
		conv1_result[5][10][4] <= 18'd0;\
		conv1_result[5][10][5] <= 18'd0;\
		conv1_result[5][10][6] <= 18'd0;\
		conv1_result[5][10][7] <= 18'd0;\
		conv1_result[5][10][8] <= 18'd0;\
		conv1_result[5][10][9] <= 18'd0;\
		conv1_result[5][10][10] <= 18'd0;\
		conv1_result[5][10][11] <= 18'd0;\
		conv1_result[5][10][12] <= 18'd0;\
		conv1_result[5][10][13] <= 18'd0;\
		conv1_result[5][11][0] <= 18'd0;\
		conv1_result[5][11][1] <= 18'd0;\
		conv1_result[5][11][2] <= 18'd0;\
		conv1_result[5][11][3] <= 18'd0;\
		conv1_result[5][11][4] <= 18'd0;\
		conv1_result[5][11][5] <= 18'd0;\
		conv1_result[5][11][6] <= 18'd0;\
		conv1_result[5][11][7] <= 18'd0;\
		conv1_result[5][11][8] <= 18'd0;\
		conv1_result[5][11][9] <= 18'd0;\
		conv1_result[5][11][10] <= 18'd0;\
		conv1_result[5][11][11] <= 18'd0;\
		conv1_result[5][11][12] <= 18'd0;\
		conv1_result[5][11][13] <= 18'd0;\
		conv1_result[5][12][0] <= 18'd0;\
		conv1_result[5][12][1] <= 18'd0;\
		conv1_result[5][12][2] <= 18'd0;\
		conv1_result[5][12][3] <= 18'd0;\
		conv1_result[5][12][4] <= 18'd0;\
		conv1_result[5][12][5] <= 18'd0;\
		conv1_result[5][12][6] <= 18'd0;\
		conv1_result[5][12][7] <= 18'd0;\
		conv1_result[5][12][8] <= 18'd0;\
		conv1_result[5][12][9] <= 18'd0;\
		conv1_result[5][12][10] <= 18'd0;\
		conv1_result[5][12][11] <= 18'd0;\
		conv1_result[5][12][12] <= 18'd0;\
		conv1_result[5][12][13] <= 18'd0;\
		conv1_result[5][13][0] <= 18'd0;\
		conv1_result[5][13][1] <= 18'd0;\
		conv1_result[5][13][2] <= 18'd0;\
		conv1_result[5][13][3] <= 18'd0;\
		conv1_result[5][13][4] <= 18'd0;\
		conv1_result[5][13][5] <= 18'd0;\
		conv1_result[5][13][6] <= 18'd0;\
		conv1_result[5][13][7] <= 18'd0;\
		conv1_result[5][13][8] <= 18'd0;\
		conv1_result[5][13][9] <= 18'd0;\
		conv1_result[5][13][10] <= 18'd0;\
		conv1_result[5][13][11] <= 18'd0;\
		conv1_result[5][13][12] <= 18'd0;\
		conv1_result[5][13][13] <= 18'd0;\
    end\
    else begin\
        case(state)\
            IDLE     :begin\
                conv1_result[0][0][0] <= 18'd0;\
                conv1_result[0][0][1] <= 18'd0;\
                conv1_result[0][0][2] <= 18'd0;\
                conv1_result[0][0][3] <= 18'd0;\
                conv1_result[0][0][4] <= 18'd0;\
                conv1_result[0][0][5] <= 18'd0;\
                conv1_result[0][0][6] <= 18'd0;\
                conv1_result[0][0][7] <= 18'd0;\
                conv1_result[0][0][8] <= 18'd0;\
                conv1_result[0][0][9] <= 18'd0;\
                conv1_result[0][0][10] <= 18'd0;\
                conv1_result[0][0][11] <= 18'd0;\
                conv1_result[0][0][12] <= 18'd0;\
                conv1_result[0][0][13] <= 18'd0;\
                conv1_result[0][1][0] <= 18'd0;\
                conv1_result[0][1][1] <= 18'd0;\
                conv1_result[0][1][2] <= 18'd0;\
                conv1_result[0][1][3] <= 18'd0;\
                conv1_result[0][1][4] <= 18'd0;\
                conv1_result[0][1][5] <= 18'd0;\
                conv1_result[0][1][6] <= 18'd0;\
                conv1_result[0][1][7] <= 18'd0;\
                conv1_result[0][1][8] <= 18'd0;\
                conv1_result[0][1][9] <= 18'd0;\
                conv1_result[0][1][10] <= 18'd0;\
                conv1_result[0][1][11] <= 18'd0;\
                conv1_result[0][1][12] <= 18'd0;\
                conv1_result[0][1][13] <= 18'd0;\
                conv1_result[0][2][0] <= 18'd0;\
                conv1_result[0][2][1] <= 18'd0;\
                conv1_result[0][2][2] <= 18'd0;\
                conv1_result[0][2][3] <= 18'd0;\
                conv1_result[0][2][4] <= 18'd0;\
                conv1_result[0][2][5] <= 18'd0;\
                conv1_result[0][2][6] <= 18'd0;\
                conv1_result[0][2][7] <= 18'd0;\
                conv1_result[0][2][8] <= 18'd0;\
                conv1_result[0][2][9] <= 18'd0;\
                conv1_result[0][2][10] <= 18'd0;\
                conv1_result[0][2][11] <= 18'd0;\
                conv1_result[0][2][12] <= 18'd0;\
                conv1_result[0][2][13] <= 18'd0;\
                conv1_result[0][3][0] <= 18'd0;\
                conv1_result[0][3][1] <= 18'd0;\
                conv1_result[0][3][2] <= 18'd0;\
                conv1_result[0][3][3] <= 18'd0;\
                conv1_result[0][3][4] <= 18'd0;\
                conv1_result[0][3][5] <= 18'd0;\
                conv1_result[0][3][6] <= 18'd0;\
                conv1_result[0][3][7] <= 18'd0;\
                conv1_result[0][3][8] <= 18'd0;\
                conv1_result[0][3][9] <= 18'd0;\
                conv1_result[0][3][10] <= 18'd0;\
                conv1_result[0][3][11] <= 18'd0;\
                conv1_result[0][3][12] <= 18'd0;\
                conv1_result[0][3][13] <= 18'd0;\
                conv1_result[0][4][0] <= 18'd0;\
                conv1_result[0][4][1] <= 18'd0;\
                conv1_result[0][4][2] <= 18'd0;\
                conv1_result[0][4][3] <= 18'd0;\
                conv1_result[0][4][4] <= 18'd0;\
                conv1_result[0][4][5] <= 18'd0;\
                conv1_result[0][4][6] <= 18'd0;\
                conv1_result[0][4][7] <= 18'd0;\
                conv1_result[0][4][8] <= 18'd0;\
                conv1_result[0][4][9] <= 18'd0;\
                conv1_result[0][4][10] <= 18'd0;\
                conv1_result[0][4][11] <= 18'd0;\
                conv1_result[0][4][12] <= 18'd0;\
                conv1_result[0][4][13] <= 18'd0;\
                conv1_result[0][5][0] <= 18'd0;\
                conv1_result[0][5][1] <= 18'd0;\
                conv1_result[0][5][2] <= 18'd0;\
                conv1_result[0][5][3] <= 18'd0;\
                conv1_result[0][5][4] <= 18'd0;\
                conv1_result[0][5][5] <= 18'd0;\
                conv1_result[0][5][6] <= 18'd0;\
                conv1_result[0][5][7] <= 18'd0;\
                conv1_result[0][5][8] <= 18'd0;\
                conv1_result[0][5][9] <= 18'd0;\
                conv1_result[0][5][10] <= 18'd0;\
                conv1_result[0][5][11] <= 18'd0;\
                conv1_result[0][5][12] <= 18'd0;\
                conv1_result[0][5][13] <= 18'd0;\
                conv1_result[0][6][0] <= 18'd0;\
                conv1_result[0][6][1] <= 18'd0;\
                conv1_result[0][6][2] <= 18'd0;\
                conv1_result[0][6][3] <= 18'd0;\
                conv1_result[0][6][4] <= 18'd0;\
                conv1_result[0][6][5] <= 18'd0;\
                conv1_result[0][6][6] <= 18'd0;\
                conv1_result[0][6][7] <= 18'd0;\
                conv1_result[0][6][8] <= 18'd0;\
                conv1_result[0][6][9] <= 18'd0;\
                conv1_result[0][6][10] <= 18'd0;\
                conv1_result[0][6][11] <= 18'd0;\
                conv1_result[0][6][12] <= 18'd0;\
                conv1_result[0][6][13] <= 18'd0;\
                conv1_result[0][7][0] <= 18'd0;\
                conv1_result[0][7][1] <= 18'd0;\
                conv1_result[0][7][2] <= 18'd0;\
                conv1_result[0][7][3] <= 18'd0;\
                conv1_result[0][7][4] <= 18'd0;\
                conv1_result[0][7][5] <= 18'd0;\
                conv1_result[0][7][6] <= 18'd0;\
                conv1_result[0][7][7] <= 18'd0;\
                conv1_result[0][7][8] <= 18'd0;\
                conv1_result[0][7][9] <= 18'd0;\
                conv1_result[0][7][10] <= 18'd0;\
                conv1_result[0][7][11] <= 18'd0;\
                conv1_result[0][7][12] <= 18'd0;\
                conv1_result[0][7][13] <= 18'd0;\
                conv1_result[0][8][0] <= 18'd0;\
                conv1_result[0][8][1] <= 18'd0;\
                conv1_result[0][8][2] <= 18'd0;\
                conv1_result[0][8][3] <= 18'd0;\
                conv1_result[0][8][4] <= 18'd0;\
                conv1_result[0][8][5] <= 18'd0;\
                conv1_result[0][8][6] <= 18'd0;\
                conv1_result[0][8][7] <= 18'd0;\
                conv1_result[0][8][8] <= 18'd0;\
                conv1_result[0][8][9] <= 18'd0;\
                conv1_result[0][8][10] <= 18'd0;\
                conv1_result[0][8][11] <= 18'd0;\
                conv1_result[0][8][12] <= 18'd0;\
                conv1_result[0][8][13] <= 18'd0;\
                conv1_result[0][9][0] <= 18'd0;\
                conv1_result[0][9][1] <= 18'd0;\
                conv1_result[0][9][2] <= 18'd0;\
                conv1_result[0][9][3] <= 18'd0;\
                conv1_result[0][9][4] <= 18'd0;\
                conv1_result[0][9][5] <= 18'd0;\
                conv1_result[0][9][6] <= 18'd0;\
                conv1_result[0][9][7] <= 18'd0;\
                conv1_result[0][9][8] <= 18'd0;\
                conv1_result[0][9][9] <= 18'd0;\
                conv1_result[0][9][10] <= 18'd0;\
                conv1_result[0][9][11] <= 18'd0;\
                conv1_result[0][9][12] <= 18'd0;\
                conv1_result[0][9][13] <= 18'd0;\
                conv1_result[0][10][0] <= 18'd0;\
                conv1_result[0][10][1] <= 18'd0;\
                conv1_result[0][10][2] <= 18'd0;\
                conv1_result[0][10][3] <= 18'd0;\
                conv1_result[0][10][4] <= 18'd0;\
                conv1_result[0][10][5] <= 18'd0;\
                conv1_result[0][10][6] <= 18'd0;\
                conv1_result[0][10][7] <= 18'd0;\
                conv1_result[0][10][8] <= 18'd0;\
                conv1_result[0][10][9] <= 18'd0;\
                conv1_result[0][10][10] <= 18'd0;\
                conv1_result[0][10][11] <= 18'd0;\
                conv1_result[0][10][12] <= 18'd0;\
                conv1_result[0][10][13] <= 18'd0;\
                conv1_result[0][11][0] <= 18'd0;\
                conv1_result[0][11][1] <= 18'd0;\
                conv1_result[0][11][2] <= 18'd0;\
                conv1_result[0][11][3] <= 18'd0;\
                conv1_result[0][11][4] <= 18'd0;\
                conv1_result[0][11][5] <= 18'd0;\
                conv1_result[0][11][6] <= 18'd0;\
                conv1_result[0][11][7] <= 18'd0;\
                conv1_result[0][11][8] <= 18'd0;\
                conv1_result[0][11][9] <= 18'd0;\
                conv1_result[0][11][10] <= 18'd0;\
                conv1_result[0][11][11] <= 18'd0;\
                conv1_result[0][11][12] <= 18'd0;\
                conv1_result[0][11][13] <= 18'd0;\
                conv1_result[0][12][0] <= 18'd0;\
                conv1_result[0][12][1] <= 18'd0;\
                conv1_result[0][12][2] <= 18'd0;\
                conv1_result[0][12][3] <= 18'd0;\
                conv1_result[0][12][4] <= 18'd0;\
                conv1_result[0][12][5] <= 18'd0;\
                conv1_result[0][12][6] <= 18'd0;\
                conv1_result[0][12][7] <= 18'd0;\
                conv1_result[0][12][8] <= 18'd0;\
                conv1_result[0][12][9] <= 18'd0;\
                conv1_result[0][12][10] <= 18'd0;\
                conv1_result[0][12][11] <= 18'd0;\
                conv1_result[0][12][12] <= 18'd0;\
                conv1_result[0][12][13] <= 18'd0;\
                conv1_result[0][13][0] <= 18'd0;\
                conv1_result[0][13][1] <= 18'd0;\
                conv1_result[0][13][2] <= 18'd0;\
                conv1_result[0][13][3] <= 18'd0;\
                conv1_result[0][13][4] <= 18'd0;\
                conv1_result[0][13][5] <= 18'd0;\
                conv1_result[0][13][6] <= 18'd0;\
                conv1_result[0][13][7] <= 18'd0;\
                conv1_result[0][13][8] <= 18'd0;\
                conv1_result[0][13][9] <= 18'd0;\
                conv1_result[0][13][10] <= 18'd0;\
                conv1_result[0][13][11] <= 18'd0;\
                conv1_result[0][13][12] <= 18'd0;\
                conv1_result[0][13][13] <= 18'd0;\
                conv1_result[1][0][0] <= 18'd0;\
                conv1_result[1][0][1] <= 18'd0;\
                conv1_result[1][0][2] <= 18'd0;\
                conv1_result[1][0][3] <= 18'd0;\
                conv1_result[1][0][4] <= 18'd0;\
                conv1_result[1][0][5] <= 18'd0;\
                conv1_result[1][0][6] <= 18'd0;\
                conv1_result[1][0][7] <= 18'd0;\
                conv1_result[1][0][8] <= 18'd0;\
                conv1_result[1][0][9] <= 18'd0;\
                conv1_result[1][0][10] <= 18'd0;\
                conv1_result[1][0][11] <= 18'd0;\
                conv1_result[1][0][12] <= 18'd0;\
                conv1_result[1][0][13] <= 18'd0;\
                conv1_result[1][1][0] <= 18'd0;\
                conv1_result[1][1][1] <= 18'd0;\
                conv1_result[1][1][2] <= 18'd0;\
                conv1_result[1][1][3] <= 18'd0;\
                conv1_result[1][1][4] <= 18'd0;\
                conv1_result[1][1][5] <= 18'd0;\
                conv1_result[1][1][6] <= 18'd0;\
                conv1_result[1][1][7] <= 18'd0;\
                conv1_result[1][1][8] <= 18'd0;\
                conv1_result[1][1][9] <= 18'd0;\
                conv1_result[1][1][10] <= 18'd0;\
                conv1_result[1][1][11] <= 18'd0;\
                conv1_result[1][1][12] <= 18'd0;\
                conv1_result[1][1][13] <= 18'd0;\
                conv1_result[1][2][0] <= 18'd0;\
                conv1_result[1][2][1] <= 18'd0;\
                conv1_result[1][2][2] <= 18'd0;\
                conv1_result[1][2][3] <= 18'd0;\
                conv1_result[1][2][4] <= 18'd0;\
                conv1_result[1][2][5] <= 18'd0;\
                conv1_result[1][2][6] <= 18'd0;\
                conv1_result[1][2][7] <= 18'd0;\
                conv1_result[1][2][8] <= 18'd0;\
                conv1_result[1][2][9] <= 18'd0;\
                conv1_result[1][2][10] <= 18'd0;\
                conv1_result[1][2][11] <= 18'd0;\
                conv1_result[1][2][12] <= 18'd0;\
                conv1_result[1][2][13] <= 18'd0;\
                conv1_result[1][3][0] <= 18'd0;\
                conv1_result[1][3][1] <= 18'd0;\
                conv1_result[1][3][2] <= 18'd0;\
                conv1_result[1][3][3] <= 18'd0;\
                conv1_result[1][3][4] <= 18'd0;\
                conv1_result[1][3][5] <= 18'd0;\
                conv1_result[1][3][6] <= 18'd0;\
                conv1_result[1][3][7] <= 18'd0;\
                conv1_result[1][3][8] <= 18'd0;\
                conv1_result[1][3][9] <= 18'd0;\
                conv1_result[1][3][10] <= 18'd0;\
                conv1_result[1][3][11] <= 18'd0;\
                conv1_result[1][3][12] <= 18'd0;\
                conv1_result[1][3][13] <= 18'd0;\
                conv1_result[1][4][0] <= 18'd0;\
                conv1_result[1][4][1] <= 18'd0;\
                conv1_result[1][4][2] <= 18'd0;\
                conv1_result[1][4][3] <= 18'd0;\
                conv1_result[1][4][4] <= 18'd0;\
                conv1_result[1][4][5] <= 18'd0;\
                conv1_result[1][4][6] <= 18'd0;\
                conv1_result[1][4][7] <= 18'd0;\
                conv1_result[1][4][8] <= 18'd0;\
                conv1_result[1][4][9] <= 18'd0;\
                conv1_result[1][4][10] <= 18'd0;\
                conv1_result[1][4][11] <= 18'd0;\
                conv1_result[1][4][12] <= 18'd0;\
                conv1_result[1][4][13] <= 18'd0;\
                conv1_result[1][5][0] <= 18'd0;\
                conv1_result[1][5][1] <= 18'd0;\
                conv1_result[1][5][2] <= 18'd0;\
                conv1_result[1][5][3] <= 18'd0;\
                conv1_result[1][5][4] <= 18'd0;\
                conv1_result[1][5][5] <= 18'd0;\
                conv1_result[1][5][6] <= 18'd0;\
                conv1_result[1][5][7] <= 18'd0;\
                conv1_result[1][5][8] <= 18'd0;\
                conv1_result[1][5][9] <= 18'd0;\
                conv1_result[1][5][10] <= 18'd0;\
                conv1_result[1][5][11] <= 18'd0;\
                conv1_result[1][5][12] <= 18'd0;\
                conv1_result[1][5][13] <= 18'd0;\
                conv1_result[1][6][0] <= 18'd0;\
                conv1_result[1][6][1] <= 18'd0;\
                conv1_result[1][6][2] <= 18'd0;\
                conv1_result[1][6][3] <= 18'd0;\
                conv1_result[1][6][4] <= 18'd0;\
                conv1_result[1][6][5] <= 18'd0;\
                conv1_result[1][6][6] <= 18'd0;\
                conv1_result[1][6][7] <= 18'd0;\
                conv1_result[1][6][8] <= 18'd0;\
                conv1_result[1][6][9] <= 18'd0;\
                conv1_result[1][6][10] <= 18'd0;\
                conv1_result[1][6][11] <= 18'd0;\
                conv1_result[1][6][12] <= 18'd0;\
                conv1_result[1][6][13] <= 18'd0;\
                conv1_result[1][7][0] <= 18'd0;\
                conv1_result[1][7][1] <= 18'd0;\
                conv1_result[1][7][2] <= 18'd0;\
                conv1_result[1][7][3] <= 18'd0;\
                conv1_result[1][7][4] <= 18'd0;\
                conv1_result[1][7][5] <= 18'd0;\
                conv1_result[1][7][6] <= 18'd0;\
                conv1_result[1][7][7] <= 18'd0;\
                conv1_result[1][7][8] <= 18'd0;\
                conv1_result[1][7][9] <= 18'd0;\
                conv1_result[1][7][10] <= 18'd0;\
                conv1_result[1][7][11] <= 18'd0;\
                conv1_result[1][7][12] <= 18'd0;\
                conv1_result[1][7][13] <= 18'd0;\
                conv1_result[1][8][0] <= 18'd0;\
                conv1_result[1][8][1] <= 18'd0;\
                conv1_result[1][8][2] <= 18'd0;\
                conv1_result[1][8][3] <= 18'd0;\
                conv1_result[1][8][4] <= 18'd0;\
                conv1_result[1][8][5] <= 18'd0;\
                conv1_result[1][8][6] <= 18'd0;\
                conv1_result[1][8][7] <= 18'd0;\
                conv1_result[1][8][8] <= 18'd0;\
                conv1_result[1][8][9] <= 18'd0;\
                conv1_result[1][8][10] <= 18'd0;\
                conv1_result[1][8][11] <= 18'd0;\
                conv1_result[1][8][12] <= 18'd0;\
                conv1_result[1][8][13] <= 18'd0;\
                conv1_result[1][9][0] <= 18'd0;\
                conv1_result[1][9][1] <= 18'd0;\
                conv1_result[1][9][2] <= 18'd0;\
                conv1_result[1][9][3] <= 18'd0;\
                conv1_result[1][9][4] <= 18'd0;\
                conv1_result[1][9][5] <= 18'd0;\
                conv1_result[1][9][6] <= 18'd0;\
                conv1_result[1][9][7] <= 18'd0;\
                conv1_result[1][9][8] <= 18'd0;\
                conv1_result[1][9][9] <= 18'd0;\
                conv1_result[1][9][10] <= 18'd0;\
                conv1_result[1][9][11] <= 18'd0;\
                conv1_result[1][9][12] <= 18'd0;\
                conv1_result[1][9][13] <= 18'd0;\
                conv1_result[1][10][0] <= 18'd0;\
                conv1_result[1][10][1] <= 18'd0;\
                conv1_result[1][10][2] <= 18'd0;\
                conv1_result[1][10][3] <= 18'd0;\
                conv1_result[1][10][4] <= 18'd0;\
                conv1_result[1][10][5] <= 18'd0;\
                conv1_result[1][10][6] <= 18'd0;\
                conv1_result[1][10][7] <= 18'd0;\
                conv1_result[1][10][8] <= 18'd0;\
                conv1_result[1][10][9] <= 18'd0;\
                conv1_result[1][10][10] <= 18'd0;\
                conv1_result[1][10][11] <= 18'd0;\
                conv1_result[1][10][12] <= 18'd0;\
                conv1_result[1][10][13] <= 18'd0;\
                conv1_result[1][11][0] <= 18'd0;\
                conv1_result[1][11][1] <= 18'd0;\
                conv1_result[1][11][2] <= 18'd0;\
                conv1_result[1][11][3] <= 18'd0;\
                conv1_result[1][11][4] <= 18'd0;\
                conv1_result[1][11][5] <= 18'd0;\
                conv1_result[1][11][6] <= 18'd0;\
                conv1_result[1][11][7] <= 18'd0;\
                conv1_result[1][11][8] <= 18'd0;\
                conv1_result[1][11][9] <= 18'd0;\
                conv1_result[1][11][10] <= 18'd0;\
                conv1_result[1][11][11] <= 18'd0;\
                conv1_result[1][11][12] <= 18'd0;\
                conv1_result[1][11][13] <= 18'd0;\
                conv1_result[1][12][0] <= 18'd0;\
                conv1_result[1][12][1] <= 18'd0;\
                conv1_result[1][12][2] <= 18'd0;\
                conv1_result[1][12][3] <= 18'd0;\
                conv1_result[1][12][4] <= 18'd0;\
                conv1_result[1][12][5] <= 18'd0;\
                conv1_result[1][12][6] <= 18'd0;\
                conv1_result[1][12][7] <= 18'd0;\
                conv1_result[1][12][8] <= 18'd0;\
                conv1_result[1][12][9] <= 18'd0;\
                conv1_result[1][12][10] <= 18'd0;\
                conv1_result[1][12][11] <= 18'd0;\
                conv1_result[1][12][12] <= 18'd0;\
                conv1_result[1][12][13] <= 18'd0;\
                conv1_result[1][13][0] <= 18'd0;\
                conv1_result[1][13][1] <= 18'd0;\
                conv1_result[1][13][2] <= 18'd0;\
                conv1_result[1][13][3] <= 18'd0;\
                conv1_result[1][13][4] <= 18'd0;\
                conv1_result[1][13][5] <= 18'd0;\
                conv1_result[1][13][6] <= 18'd0;\
                conv1_result[1][13][7] <= 18'd0;\
                conv1_result[1][13][8] <= 18'd0;\
                conv1_result[1][13][9] <= 18'd0;\
                conv1_result[1][13][10] <= 18'd0;\
                conv1_result[1][13][11] <= 18'd0;\
                conv1_result[1][13][12] <= 18'd0;\
                conv1_result[1][13][13] <= 18'd0;\
                conv1_result[2][0][0] <= 18'd0;\
                conv1_result[2][0][1] <= 18'd0;\
                conv1_result[2][0][2] <= 18'd0;\
                conv1_result[2][0][3] <= 18'd0;\
                conv1_result[2][0][4] <= 18'd0;\
                conv1_result[2][0][5] <= 18'd0;\
                conv1_result[2][0][6] <= 18'd0;\
                conv1_result[2][0][7] <= 18'd0;\
                conv1_result[2][0][8] <= 18'd0;\
                conv1_result[2][0][9] <= 18'd0;\
                conv1_result[2][0][10] <= 18'd0;\
                conv1_result[2][0][11] <= 18'd0;\
                conv1_result[2][0][12] <= 18'd0;\
                conv1_result[2][0][13] <= 18'd0;\
                conv1_result[2][1][0] <= 18'd0;\
                conv1_result[2][1][1] <= 18'd0;\
                conv1_result[2][1][2] <= 18'd0;\
                conv1_result[2][1][3] <= 18'd0;\
                conv1_result[2][1][4] <= 18'd0;\
                conv1_result[2][1][5] <= 18'd0;\
                conv1_result[2][1][6] <= 18'd0;\
                conv1_result[2][1][7] <= 18'd0;\
                conv1_result[2][1][8] <= 18'd0;\
                conv1_result[2][1][9] <= 18'd0;\
                conv1_result[2][1][10] <= 18'd0;\
                conv1_result[2][1][11] <= 18'd0;\
                conv1_result[2][1][12] <= 18'd0;\
                conv1_result[2][1][13] <= 18'd0;\
                conv1_result[2][2][0] <= 18'd0;\
                conv1_result[2][2][1] <= 18'd0;\
                conv1_result[2][2][2] <= 18'd0;\
                conv1_result[2][2][3] <= 18'd0;\
                conv1_result[2][2][4] <= 18'd0;\
                conv1_result[2][2][5] <= 18'd0;\
                conv1_result[2][2][6] <= 18'd0;\
                conv1_result[2][2][7] <= 18'd0;\
                conv1_result[2][2][8] <= 18'd0;\
                conv1_result[2][2][9] <= 18'd0;\
                conv1_result[2][2][10] <= 18'd0;\
                conv1_result[2][2][11] <= 18'd0;\
                conv1_result[2][2][12] <= 18'd0;\
                conv1_result[2][2][13] <= 18'd0;\
                conv1_result[2][3][0] <= 18'd0;\
                conv1_result[2][3][1] <= 18'd0;\
                conv1_result[2][3][2] <= 18'd0;\
                conv1_result[2][3][3] <= 18'd0;\
                conv1_result[2][3][4] <= 18'd0;\
                conv1_result[2][3][5] <= 18'd0;\
                conv1_result[2][3][6] <= 18'd0;\
                conv1_result[2][3][7] <= 18'd0;\
                conv1_result[2][3][8] <= 18'd0;\
                conv1_result[2][3][9] <= 18'd0;\
                conv1_result[2][3][10] <= 18'd0;\
                conv1_result[2][3][11] <= 18'd0;\
                conv1_result[2][3][12] <= 18'd0;\
                conv1_result[2][3][13] <= 18'd0;\
                conv1_result[2][4][0] <= 18'd0;\
                conv1_result[2][4][1] <= 18'd0;\
                conv1_result[2][4][2] <= 18'd0;\
                conv1_result[2][4][3] <= 18'd0;\
                conv1_result[2][4][4] <= 18'd0;\
                conv1_result[2][4][5] <= 18'd0;\
                conv1_result[2][4][6] <= 18'd0;\
                conv1_result[2][4][7] <= 18'd0;\
                conv1_result[2][4][8] <= 18'd0;\
                conv1_result[2][4][9] <= 18'd0;\
                conv1_result[2][4][10] <= 18'd0;\
                conv1_result[2][4][11] <= 18'd0;\
                conv1_result[2][4][12] <= 18'd0;\
                conv1_result[2][4][13] <= 18'd0;\
                conv1_result[2][5][0] <= 18'd0;\
                conv1_result[2][5][1] <= 18'd0;\
                conv1_result[2][5][2] <= 18'd0;\
                conv1_result[2][5][3] <= 18'd0;\
                conv1_result[2][5][4] <= 18'd0;\
                conv1_result[2][5][5] <= 18'd0;\
                conv1_result[2][5][6] <= 18'd0;\
                conv1_result[2][5][7] <= 18'd0;\
                conv1_result[2][5][8] <= 18'd0;\
                conv1_result[2][5][9] <= 18'd0;\
                conv1_result[2][5][10] <= 18'd0;\
                conv1_result[2][5][11] <= 18'd0;\
                conv1_result[2][5][12] <= 18'd0;\
                conv1_result[2][5][13] <= 18'd0;\
                conv1_result[2][6][0] <= 18'd0;\
                conv1_result[2][6][1] <= 18'd0;\
                conv1_result[2][6][2] <= 18'd0;\
                conv1_result[2][6][3] <= 18'd0;\
                conv1_result[2][6][4] <= 18'd0;\
                conv1_result[2][6][5] <= 18'd0;\
                conv1_result[2][6][6] <= 18'd0;\
                conv1_result[2][6][7] <= 18'd0;\
                conv1_result[2][6][8] <= 18'd0;\
                conv1_result[2][6][9] <= 18'd0;\
                conv1_result[2][6][10] <= 18'd0;\
                conv1_result[2][6][11] <= 18'd0;\
                conv1_result[2][6][12] <= 18'd0;\
                conv1_result[2][6][13] <= 18'd0;\
                conv1_result[2][7][0] <= 18'd0;\
                conv1_result[2][7][1] <= 18'd0;\
                conv1_result[2][7][2] <= 18'd0;\
                conv1_result[2][7][3] <= 18'd0;\
                conv1_result[2][7][4] <= 18'd0;\
                conv1_result[2][7][5] <= 18'd0;\
                conv1_result[2][7][6] <= 18'd0;\
                conv1_result[2][7][7] <= 18'd0;\
                conv1_result[2][7][8] <= 18'd0;\
                conv1_result[2][7][9] <= 18'd0;\
                conv1_result[2][7][10] <= 18'd0;\
                conv1_result[2][7][11] <= 18'd0;\
                conv1_result[2][7][12] <= 18'd0;\
                conv1_result[2][7][13] <= 18'd0;\
                conv1_result[2][8][0] <= 18'd0;\
                conv1_result[2][8][1] <= 18'd0;\
                conv1_result[2][8][2] <= 18'd0;\
                conv1_result[2][8][3] <= 18'd0;\
                conv1_result[2][8][4] <= 18'd0;\
                conv1_result[2][8][5] <= 18'd0;\
                conv1_result[2][8][6] <= 18'd0;\
                conv1_result[2][8][7] <= 18'd0;\
                conv1_result[2][8][8] <= 18'd0;\
                conv1_result[2][8][9] <= 18'd0;\
                conv1_result[2][8][10] <= 18'd0;\
                conv1_result[2][8][11] <= 18'd0;\
                conv1_result[2][8][12] <= 18'd0;\
                conv1_result[2][8][13] <= 18'd0;\
                conv1_result[2][9][0] <= 18'd0;\
                conv1_result[2][9][1] <= 18'd0;\
                conv1_result[2][9][2] <= 18'd0;\
                conv1_result[2][9][3] <= 18'd0;\
                conv1_result[2][9][4] <= 18'd0;\
                conv1_result[2][9][5] <= 18'd0;\
                conv1_result[2][9][6] <= 18'd0;\
                conv1_result[2][9][7] <= 18'd0;\
                conv1_result[2][9][8] <= 18'd0;\
                conv1_result[2][9][9] <= 18'd0;\
                conv1_result[2][9][10] <= 18'd0;\
                conv1_result[2][9][11] <= 18'd0;\
                conv1_result[2][9][12] <= 18'd0;\
                conv1_result[2][9][13] <= 18'd0;\
                conv1_result[2][10][0] <= 18'd0;\
                conv1_result[2][10][1] <= 18'd0;\
                conv1_result[2][10][2] <= 18'd0;\
                conv1_result[2][10][3] <= 18'd0;\
                conv1_result[2][10][4] <= 18'd0;\
                conv1_result[2][10][5] <= 18'd0;\
                conv1_result[2][10][6] <= 18'd0;\
                conv1_result[2][10][7] <= 18'd0;\
                conv1_result[2][10][8] <= 18'd0;\
                conv1_result[2][10][9] <= 18'd0;\
                conv1_result[2][10][10] <= 18'd0;\
                conv1_result[2][10][11] <= 18'd0;\
                conv1_result[2][10][12] <= 18'd0;\
                conv1_result[2][10][13] <= 18'd0;\
                conv1_result[2][11][0] <= 18'd0;\
                conv1_result[2][11][1] <= 18'd0;\
                conv1_result[2][11][2] <= 18'd0;\
                conv1_result[2][11][3] <= 18'd0;\
                conv1_result[2][11][4] <= 18'd0;\
                conv1_result[2][11][5] <= 18'd0;\
                conv1_result[2][11][6] <= 18'd0;\
                conv1_result[2][11][7] <= 18'd0;\
                conv1_result[2][11][8] <= 18'd0;\
                conv1_result[2][11][9] <= 18'd0;\
                conv1_result[2][11][10] <= 18'd0;\
                conv1_result[2][11][11] <= 18'd0;\
                conv1_result[2][11][12] <= 18'd0;\
                conv1_result[2][11][13] <= 18'd0;\
                conv1_result[2][12][0] <= 18'd0;\
                conv1_result[2][12][1] <= 18'd0;\
                conv1_result[2][12][2] <= 18'd0;\
                conv1_result[2][12][3] <= 18'd0;\
                conv1_result[2][12][4] <= 18'd0;\
                conv1_result[2][12][5] <= 18'd0;\
                conv1_result[2][12][6] <= 18'd0;\
                conv1_result[2][12][7] <= 18'd0;\
                conv1_result[2][12][8] <= 18'd0;\
                conv1_result[2][12][9] <= 18'd0;\
                conv1_result[2][12][10] <= 18'd0;\
                conv1_result[2][12][11] <= 18'd0;\
                conv1_result[2][12][12] <= 18'd0;\
                conv1_result[2][12][13] <= 18'd0;\
                conv1_result[2][13][0] <= 18'd0;\
                conv1_result[2][13][1] <= 18'd0;\
                conv1_result[2][13][2] <= 18'd0;\
                conv1_result[2][13][3] <= 18'd0;\
                conv1_result[2][13][4] <= 18'd0;\
                conv1_result[2][13][5] <= 18'd0;\
                conv1_result[2][13][6] <= 18'd0;\
                conv1_result[2][13][7] <= 18'd0;\
                conv1_result[2][13][8] <= 18'd0;\
                conv1_result[2][13][9] <= 18'd0;\
                conv1_result[2][13][10] <= 18'd0;\
                conv1_result[2][13][11] <= 18'd0;\
                conv1_result[2][13][12] <= 18'd0;\
                conv1_result[2][13][13] <= 18'd0;\
                conv1_result[3][0][0] <= 18'd0;\
                conv1_result[3][0][1] <= 18'd0;\
                conv1_result[3][0][2] <= 18'd0;\
                conv1_result[3][0][3] <= 18'd0;\
                conv1_result[3][0][4] <= 18'd0;\
                conv1_result[3][0][5] <= 18'd0;\
                conv1_result[3][0][6] <= 18'd0;\
                conv1_result[3][0][7] <= 18'd0;\
                conv1_result[3][0][8] <= 18'd0;\
                conv1_result[3][0][9] <= 18'd0;\
                conv1_result[3][0][10] <= 18'd0;\
                conv1_result[3][0][11] <= 18'd0;\
                conv1_result[3][0][12] <= 18'd0;\
                conv1_result[3][0][13] <= 18'd0;\
                conv1_result[3][1][0] <= 18'd0;\
                conv1_result[3][1][1] <= 18'd0;\
                conv1_result[3][1][2] <= 18'd0;\
                conv1_result[3][1][3] <= 18'd0;\
                conv1_result[3][1][4] <= 18'd0;\
                conv1_result[3][1][5] <= 18'd0;\
                conv1_result[3][1][6] <= 18'd0;\
                conv1_result[3][1][7] <= 18'd0;\
                conv1_result[3][1][8] <= 18'd0;\
                conv1_result[3][1][9] <= 18'd0;\
                conv1_result[3][1][10] <= 18'd0;\
                conv1_result[3][1][11] <= 18'd0;\
                conv1_result[3][1][12] <= 18'd0;\
                conv1_result[3][1][13] <= 18'd0;\
                conv1_result[3][2][0] <= 18'd0;\
                conv1_result[3][2][1] <= 18'd0;\
                conv1_result[3][2][2] <= 18'd0;\
                conv1_result[3][2][3] <= 18'd0;\
                conv1_result[3][2][4] <= 18'd0;\
                conv1_result[3][2][5] <= 18'd0;\
                conv1_result[3][2][6] <= 18'd0;\
                conv1_result[3][2][7] <= 18'd0;\
                conv1_result[3][2][8] <= 18'd0;\
                conv1_result[3][2][9] <= 18'd0;\
                conv1_result[3][2][10] <= 18'd0;\
                conv1_result[3][2][11] <= 18'd0;\
                conv1_result[3][2][12] <= 18'd0;\
                conv1_result[3][2][13] <= 18'd0;\
                conv1_result[3][3][0] <= 18'd0;\
                conv1_result[3][3][1] <= 18'd0;\
                conv1_result[3][3][2] <= 18'd0;\
                conv1_result[3][3][3] <= 18'd0;\
                conv1_result[3][3][4] <= 18'd0;\
                conv1_result[3][3][5] <= 18'd0;\
                conv1_result[3][3][6] <= 18'd0;\
                conv1_result[3][3][7] <= 18'd0;\
                conv1_result[3][3][8] <= 18'd0;\
                conv1_result[3][3][9] <= 18'd0;\
                conv1_result[3][3][10] <= 18'd0;\
                conv1_result[3][3][11] <= 18'd0;\
                conv1_result[3][3][12] <= 18'd0;\
                conv1_result[3][3][13] <= 18'd0;\
                conv1_result[3][4][0] <= 18'd0;\
                conv1_result[3][4][1] <= 18'd0;\
                conv1_result[3][4][2] <= 18'd0;\
                conv1_result[3][4][3] <= 18'd0;\
                conv1_result[3][4][4] <= 18'd0;\
                conv1_result[3][4][5] <= 18'd0;\
                conv1_result[3][4][6] <= 18'd0;\
                conv1_result[3][4][7] <= 18'd0;\
                conv1_result[3][4][8] <= 18'd0;\
                conv1_result[3][4][9] <= 18'd0;\
                conv1_result[3][4][10] <= 18'd0;\
                conv1_result[3][4][11] <= 18'd0;\
                conv1_result[3][4][12] <= 18'd0;\
                conv1_result[3][4][13] <= 18'd0;\
                conv1_result[3][5][0] <= 18'd0;\
                conv1_result[3][5][1] <= 18'd0;\
                conv1_result[3][5][2] <= 18'd0;\
                conv1_result[3][5][3] <= 18'd0;\
                conv1_result[3][5][4] <= 18'd0;\
                conv1_result[3][5][5] <= 18'd0;\
                conv1_result[3][5][6] <= 18'd0;\
                conv1_result[3][5][7] <= 18'd0;\
                conv1_result[3][5][8] <= 18'd0;\
                conv1_result[3][5][9] <= 18'd0;\
                conv1_result[3][5][10] <= 18'd0;\
                conv1_result[3][5][11] <= 18'd0;\
                conv1_result[3][5][12] <= 18'd0;\
                conv1_result[3][5][13] <= 18'd0;\
                conv1_result[3][6][0] <= 18'd0;\
                conv1_result[3][6][1] <= 18'd0;\
                conv1_result[3][6][2] <= 18'd0;\
                conv1_result[3][6][3] <= 18'd0;\
                conv1_result[3][6][4] <= 18'd0;\
                conv1_result[3][6][5] <= 18'd0;\
                conv1_result[3][6][6] <= 18'd0;\
                conv1_result[3][6][7] <= 18'd0;\
                conv1_result[3][6][8] <= 18'd0;\
                conv1_result[3][6][9] <= 18'd0;\
                conv1_result[3][6][10] <= 18'd0;\
                conv1_result[3][6][11] <= 18'd0;\
                conv1_result[3][6][12] <= 18'd0;\
                conv1_result[3][6][13] <= 18'd0;\
                conv1_result[3][7][0] <= 18'd0;\
                conv1_result[3][7][1] <= 18'd0;\
                conv1_result[3][7][2] <= 18'd0;\
                conv1_result[3][7][3] <= 18'd0;\
                conv1_result[3][7][4] <= 18'd0;\
                conv1_result[3][7][5] <= 18'd0;\
                conv1_result[3][7][6] <= 18'd0;\
                conv1_result[3][7][7] <= 18'd0;\
                conv1_result[3][7][8] <= 18'd0;\
                conv1_result[3][7][9] <= 18'd0;\
                conv1_result[3][7][10] <= 18'd0;\
                conv1_result[3][7][11] <= 18'd0;\
                conv1_result[3][7][12] <= 18'd0;\
                conv1_result[3][7][13] <= 18'd0;\
                conv1_result[3][8][0] <= 18'd0;\
                conv1_result[3][8][1] <= 18'd0;\
                conv1_result[3][8][2] <= 18'd0;\
                conv1_result[3][8][3] <= 18'd0;\
                conv1_result[3][8][4] <= 18'd0;\
                conv1_result[3][8][5] <= 18'd0;\
                conv1_result[3][8][6] <= 18'd0;\
                conv1_result[3][8][7] <= 18'd0;\
                conv1_result[3][8][8] <= 18'd0;\
                conv1_result[3][8][9] <= 18'd0;\
                conv1_result[3][8][10] <= 18'd0;\
                conv1_result[3][8][11] <= 18'd0;\
                conv1_result[3][8][12] <= 18'd0;\
                conv1_result[3][8][13] <= 18'd0;\
                conv1_result[3][9][0] <= 18'd0;\
                conv1_result[3][9][1] <= 18'd0;\
                conv1_result[3][9][2] <= 18'd0;\
                conv1_result[3][9][3] <= 18'd0;\
                conv1_result[3][9][4] <= 18'd0;\
                conv1_result[3][9][5] <= 18'd0;\
                conv1_result[3][9][6] <= 18'd0;\
                conv1_result[3][9][7] <= 18'd0;\
                conv1_result[3][9][8] <= 18'd0;\
                conv1_result[3][9][9] <= 18'd0;\
                conv1_result[3][9][10] <= 18'd0;\
                conv1_result[3][9][11] <= 18'd0;\
                conv1_result[3][9][12] <= 18'd0;\
                conv1_result[3][9][13] <= 18'd0;\
                conv1_result[3][10][0] <= 18'd0;\
                conv1_result[3][10][1] <= 18'd0;\
                conv1_result[3][10][2] <= 18'd0;\
                conv1_result[3][10][3] <= 18'd0;\
                conv1_result[3][10][4] <= 18'd0;\
                conv1_result[3][10][5] <= 18'd0;\
                conv1_result[3][10][6] <= 18'd0;\
                conv1_result[3][10][7] <= 18'd0;\
                conv1_result[3][10][8] <= 18'd0;\
                conv1_result[3][10][9] <= 18'd0;\
                conv1_result[3][10][10] <= 18'd0;\
                conv1_result[3][10][11] <= 18'd0;\
                conv1_result[3][10][12] <= 18'd0;\
                conv1_result[3][10][13] <= 18'd0;\
                conv1_result[3][11][0] <= 18'd0;\
                conv1_result[3][11][1] <= 18'd0;\
                conv1_result[3][11][2] <= 18'd0;\
                conv1_result[3][11][3] <= 18'd0;\
                conv1_result[3][11][4] <= 18'd0;\
                conv1_result[3][11][5] <= 18'd0;\
                conv1_result[3][11][6] <= 18'd0;\
                conv1_result[3][11][7] <= 18'd0;\
                conv1_result[3][11][8] <= 18'd0;\
                conv1_result[3][11][9] <= 18'd0;\
                conv1_result[3][11][10] <= 18'd0;\
                conv1_result[3][11][11] <= 18'd0;\
                conv1_result[3][11][12] <= 18'd0;\
                conv1_result[3][11][13] <= 18'd0;\
                conv1_result[3][12][0] <= 18'd0;\
                conv1_result[3][12][1] <= 18'd0;\
                conv1_result[3][12][2] <= 18'd0;\
                conv1_result[3][12][3] <= 18'd0;\
                conv1_result[3][12][4] <= 18'd0;\
                conv1_result[3][12][5] <= 18'd0;\
                conv1_result[3][12][6] <= 18'd0;\
                conv1_result[3][12][7] <= 18'd0;\
                conv1_result[3][12][8] <= 18'd0;\
                conv1_result[3][12][9] <= 18'd0;\
                conv1_result[3][12][10] <= 18'd0;\
                conv1_result[3][12][11] <= 18'd0;\
                conv1_result[3][12][12] <= 18'd0;\
                conv1_result[3][12][13] <= 18'd0;\
                conv1_result[3][13][0] <= 18'd0;\
                conv1_result[3][13][1] <= 18'd0;\
                conv1_result[3][13][2] <= 18'd0;\
                conv1_result[3][13][3] <= 18'd0;\
                conv1_result[3][13][4] <= 18'd0;\
                conv1_result[3][13][5] <= 18'd0;\
                conv1_result[3][13][6] <= 18'd0;\
                conv1_result[3][13][7] <= 18'd0;\
                conv1_result[3][13][8] <= 18'd0;\
                conv1_result[3][13][9] <= 18'd0;\
                conv1_result[3][13][10] <= 18'd0;\
                conv1_result[3][13][11] <= 18'd0;\
                conv1_result[3][13][12] <= 18'd0;\
                conv1_result[3][13][13] <= 18'd0;\
                conv1_result[4][0][0] <= 18'd0;\
                conv1_result[4][0][1] <= 18'd0;\
                conv1_result[4][0][2] <= 18'd0;\
                conv1_result[4][0][3] <= 18'd0;\
                conv1_result[4][0][4] <= 18'd0;\
                conv1_result[4][0][5] <= 18'd0;\
                conv1_result[4][0][6] <= 18'd0;\
                conv1_result[4][0][7] <= 18'd0;\
                conv1_result[4][0][8] <= 18'd0;\
                conv1_result[4][0][9] <= 18'd0;\
                conv1_result[4][0][10] <= 18'd0;\
                conv1_result[4][0][11] <= 18'd0;\
                conv1_result[4][0][12] <= 18'd0;\
                conv1_result[4][0][13] <= 18'd0;\
                conv1_result[4][1][0] <= 18'd0;\
                conv1_result[4][1][1] <= 18'd0;\
                conv1_result[4][1][2] <= 18'd0;\
                conv1_result[4][1][3] <= 18'd0;\
                conv1_result[4][1][4] <= 18'd0;\
                conv1_result[4][1][5] <= 18'd0;\
                conv1_result[4][1][6] <= 18'd0;\
                conv1_result[4][1][7] <= 18'd0;\
                conv1_result[4][1][8] <= 18'd0;\
                conv1_result[4][1][9] <= 18'd0;\
                conv1_result[4][1][10] <= 18'd0;\
                conv1_result[4][1][11] <= 18'd0;\
                conv1_result[4][1][12] <= 18'd0;\
                conv1_result[4][1][13] <= 18'd0;\
                conv1_result[4][2][0] <= 18'd0;\
                conv1_result[4][2][1] <= 18'd0;\
                conv1_result[4][2][2] <= 18'd0;\
                conv1_result[4][2][3] <= 18'd0;\
                conv1_result[4][2][4] <= 18'd0;\
                conv1_result[4][2][5] <= 18'd0;\
                conv1_result[4][2][6] <= 18'd0;\
                conv1_result[4][2][7] <= 18'd0;\
                conv1_result[4][2][8] <= 18'd0;\
                conv1_result[4][2][9] <= 18'd0;\
                conv1_result[4][2][10] <= 18'd0;\
                conv1_result[4][2][11] <= 18'd0;\
                conv1_result[4][2][12] <= 18'd0;\
                conv1_result[4][2][13] <= 18'd0;\
                conv1_result[4][3][0] <= 18'd0;\
                conv1_result[4][3][1] <= 18'd0;\
                conv1_result[4][3][2] <= 18'd0;\
                conv1_result[4][3][3] <= 18'd0;\
                conv1_result[4][3][4] <= 18'd0;\
                conv1_result[4][3][5] <= 18'd0;\
                conv1_result[4][3][6] <= 18'd0;\
                conv1_result[4][3][7] <= 18'd0;\
                conv1_result[4][3][8] <= 18'd0;\
                conv1_result[4][3][9] <= 18'd0;\
                conv1_result[4][3][10] <= 18'd0;\
                conv1_result[4][3][11] <= 18'd0;\
                conv1_result[4][3][12] <= 18'd0;\
                conv1_result[4][3][13] <= 18'd0;\
                conv1_result[4][4][0] <= 18'd0;\
                conv1_result[4][4][1] <= 18'd0;\
                conv1_result[4][4][2] <= 18'd0;\
                conv1_result[4][4][3] <= 18'd0;\
                conv1_result[4][4][4] <= 18'd0;\
                conv1_result[4][4][5] <= 18'd0;\
                conv1_result[4][4][6] <= 18'd0;\
                conv1_result[4][4][7] <= 18'd0;\
                conv1_result[4][4][8] <= 18'd0;\
                conv1_result[4][4][9] <= 18'd0;\
                conv1_result[4][4][10] <= 18'd0;\
                conv1_result[4][4][11] <= 18'd0;\
                conv1_result[4][4][12] <= 18'd0;\
                conv1_result[4][4][13] <= 18'd0;\
                conv1_result[4][5][0] <= 18'd0;\
                conv1_result[4][5][1] <= 18'd0;\
                conv1_result[4][5][2] <= 18'd0;\
                conv1_result[4][5][3] <= 18'd0;\
                conv1_result[4][5][4] <= 18'd0;\
                conv1_result[4][5][5] <= 18'd0;\
                conv1_result[4][5][6] <= 18'd0;\
                conv1_result[4][5][7] <= 18'd0;\
                conv1_result[4][5][8] <= 18'd0;\
                conv1_result[4][5][9] <= 18'd0;\
                conv1_result[4][5][10] <= 18'd0;\
                conv1_result[4][5][11] <= 18'd0;\
                conv1_result[4][5][12] <= 18'd0;\
                conv1_result[4][5][13] <= 18'd0;\
                conv1_result[4][6][0] <= 18'd0;\
                conv1_result[4][6][1] <= 18'd0;\
                conv1_result[4][6][2] <= 18'd0;\
                conv1_result[4][6][3] <= 18'd0;\
                conv1_result[4][6][4] <= 18'd0;\
                conv1_result[4][6][5] <= 18'd0;\
                conv1_result[4][6][6] <= 18'd0;\
                conv1_result[4][6][7] <= 18'd0;\
                conv1_result[4][6][8] <= 18'd0;\
                conv1_result[4][6][9] <= 18'd0;\
                conv1_result[4][6][10] <= 18'd0;\
                conv1_result[4][6][11] <= 18'd0;\
                conv1_result[4][6][12] <= 18'd0;\
                conv1_result[4][6][13] <= 18'd0;\
                conv1_result[4][7][0] <= 18'd0;\
                conv1_result[4][7][1] <= 18'd0;\
                conv1_result[4][7][2] <= 18'd0;\
                conv1_result[4][7][3] <= 18'd0;\
                conv1_result[4][7][4] <= 18'd0;\
                conv1_result[4][7][5] <= 18'd0;\
                conv1_result[4][7][6] <= 18'd0;\
                conv1_result[4][7][7] <= 18'd0;\
                conv1_result[4][7][8] <= 18'd0;\
                conv1_result[4][7][9] <= 18'd0;\
                conv1_result[4][7][10] <= 18'd0;\
                conv1_result[4][7][11] <= 18'd0;\
                conv1_result[4][7][12] <= 18'd0;\
                conv1_result[4][7][13] <= 18'd0;\
                conv1_result[4][8][0] <= 18'd0;\
                conv1_result[4][8][1] <= 18'd0;\
                conv1_result[4][8][2] <= 18'd0;\
                conv1_result[4][8][3] <= 18'd0;\
                conv1_result[4][8][4] <= 18'd0;\
                conv1_result[4][8][5] <= 18'd0;\
                conv1_result[4][8][6] <= 18'd0;\
                conv1_result[4][8][7] <= 18'd0;\
                conv1_result[4][8][8] <= 18'd0;\
                conv1_result[4][8][9] <= 18'd0;\
                conv1_result[4][8][10] <= 18'd0;\
                conv1_result[4][8][11] <= 18'd0;\
                conv1_result[4][8][12] <= 18'd0;\
                conv1_result[4][8][13] <= 18'd0;\
                conv1_result[4][9][0] <= 18'd0;\
                conv1_result[4][9][1] <= 18'd0;\
                conv1_result[4][9][2] <= 18'd0;\
                conv1_result[4][9][3] <= 18'd0;\
                conv1_result[4][9][4] <= 18'd0;\
                conv1_result[4][9][5] <= 18'd0;\
                conv1_result[4][9][6] <= 18'd0;\
                conv1_result[4][9][7] <= 18'd0;\
                conv1_result[4][9][8] <= 18'd0;\
                conv1_result[4][9][9] <= 18'd0;\
                conv1_result[4][9][10] <= 18'd0;\
                conv1_result[4][9][11] <= 18'd0;\
                conv1_result[4][9][12] <= 18'd0;\
                conv1_result[4][9][13] <= 18'd0;\
                conv1_result[4][10][0] <= 18'd0;\
                conv1_result[4][10][1] <= 18'd0;\
                conv1_result[4][10][2] <= 18'd0;\
                conv1_result[4][10][3] <= 18'd0;\
                conv1_result[4][10][4] <= 18'd0;\
                conv1_result[4][10][5] <= 18'd0;\
                conv1_result[4][10][6] <= 18'd0;\
                conv1_result[4][10][7] <= 18'd0;\
                conv1_result[4][10][8] <= 18'd0;\
                conv1_result[4][10][9] <= 18'd0;\
                conv1_result[4][10][10] <= 18'd0;\
                conv1_result[4][10][11] <= 18'd0;\
                conv1_result[4][10][12] <= 18'd0;\
                conv1_result[4][10][13] <= 18'd0;\
                conv1_result[4][11][0] <= 18'd0;\
                conv1_result[4][11][1] <= 18'd0;\
                conv1_result[4][11][2] <= 18'd0;\
                conv1_result[4][11][3] <= 18'd0;\
                conv1_result[4][11][4] <= 18'd0;\
                conv1_result[4][11][5] <= 18'd0;\
                conv1_result[4][11][6] <= 18'd0;\
                conv1_result[4][11][7] <= 18'd0;\
                conv1_result[4][11][8] <= 18'd0;\
                conv1_result[4][11][9] <= 18'd0;\
                conv1_result[4][11][10] <= 18'd0;\
                conv1_result[4][11][11] <= 18'd0;\
                conv1_result[4][11][12] <= 18'd0;\
                conv1_result[4][11][13] <= 18'd0;\
                conv1_result[4][12][0] <= 18'd0;\
                conv1_result[4][12][1] <= 18'd0;\
                conv1_result[4][12][2] <= 18'd0;\
                conv1_result[4][12][3] <= 18'd0;\
                conv1_result[4][12][4] <= 18'd0;\
                conv1_result[4][12][5] <= 18'd0;\
                conv1_result[4][12][6] <= 18'd0;\
                conv1_result[4][12][7] <= 18'd0;\
                conv1_result[4][12][8] <= 18'd0;\
                conv1_result[4][12][9] <= 18'd0;\
                conv1_result[4][12][10] <= 18'd0;\
                conv1_result[4][12][11] <= 18'd0;\
                conv1_result[4][12][12] <= 18'd0;\
                conv1_result[4][12][13] <= 18'd0;\
                conv1_result[4][13][0] <= 18'd0;\
                conv1_result[4][13][1] <= 18'd0;\
                conv1_result[4][13][2] <= 18'd0;\
                conv1_result[4][13][3] <= 18'd0;\
                conv1_result[4][13][4] <= 18'd0;\
                conv1_result[4][13][5] <= 18'd0;\
                conv1_result[4][13][6] <= 18'd0;\
                conv1_result[4][13][7] <= 18'd0;\
                conv1_result[4][13][8] <= 18'd0;\
                conv1_result[4][13][9] <= 18'd0;\
                conv1_result[4][13][10] <= 18'd0;\
                conv1_result[4][13][11] <= 18'd0;\
                conv1_result[4][13][12] <= 18'd0;\
                conv1_result[4][13][13] <= 18'd0;\
                conv1_result[5][0][0] <= 18'd0;\
                conv1_result[5][0][1] <= 18'd0;\
                conv1_result[5][0][2] <= 18'd0;\
                conv1_result[5][0][3] <= 18'd0;\
                conv1_result[5][0][4] <= 18'd0;\
                conv1_result[5][0][5] <= 18'd0;\
                conv1_result[5][0][6] <= 18'd0;\
                conv1_result[5][0][7] <= 18'd0;\
                conv1_result[5][0][8] <= 18'd0;\
                conv1_result[5][0][9] <= 18'd0;\
                conv1_result[5][0][10] <= 18'd0;\
                conv1_result[5][0][11] <= 18'd0;\
                conv1_result[5][0][12] <= 18'd0;\
                conv1_result[5][0][13] <= 18'd0;\
                conv1_result[5][1][0] <= 18'd0;\
                conv1_result[5][1][1] <= 18'd0;\
                conv1_result[5][1][2] <= 18'd0;\
                conv1_result[5][1][3] <= 18'd0;\
                conv1_result[5][1][4] <= 18'd0;\
                conv1_result[5][1][5] <= 18'd0;\
                conv1_result[5][1][6] <= 18'd0;\
                conv1_result[5][1][7] <= 18'd0;\
                conv1_result[5][1][8] <= 18'd0;\
                conv1_result[5][1][9] <= 18'd0;\
                conv1_result[5][1][10] <= 18'd0;\
                conv1_result[5][1][11] <= 18'd0;\
                conv1_result[5][1][12] <= 18'd0;\
                conv1_result[5][1][13] <= 18'd0;\
                conv1_result[5][2][0] <= 18'd0;\
                conv1_result[5][2][1] <= 18'd0;\
                conv1_result[5][2][2] <= 18'd0;\
                conv1_result[5][2][3] <= 18'd0;\
                conv1_result[5][2][4] <= 18'd0;\
                conv1_result[5][2][5] <= 18'd0;\
                conv1_result[5][2][6] <= 18'd0;\
                conv1_result[5][2][7] <= 18'd0;\
                conv1_result[5][2][8] <= 18'd0;\
                conv1_result[5][2][9] <= 18'd0;\
                conv1_result[5][2][10] <= 18'd0;\
                conv1_result[5][2][11] <= 18'd0;\
                conv1_result[5][2][12] <= 18'd0;\
                conv1_result[5][2][13] <= 18'd0;\
                conv1_result[5][3][0] <= 18'd0;\
                conv1_result[5][3][1] <= 18'd0;\
                conv1_result[5][3][2] <= 18'd0;\
                conv1_result[5][3][3] <= 18'd0;\
                conv1_result[5][3][4] <= 18'd0;\
                conv1_result[5][3][5] <= 18'd0;\
                conv1_result[5][3][6] <= 18'd0;\
                conv1_result[5][3][7] <= 18'd0;\
                conv1_result[5][3][8] <= 18'd0;\
                conv1_result[5][3][9] <= 18'd0;\
                conv1_result[5][3][10] <= 18'd0;\
                conv1_result[5][3][11] <= 18'd0;\
                conv1_result[5][3][12] <= 18'd0;\
                conv1_result[5][3][13] <= 18'd0;\
                conv1_result[5][4][0] <= 18'd0;\
                conv1_result[5][4][1] <= 18'd0;\
                conv1_result[5][4][2] <= 18'd0;\
                conv1_result[5][4][3] <= 18'd0;\
                conv1_result[5][4][4] <= 18'd0;\
                conv1_result[5][4][5] <= 18'd0;\
                conv1_result[5][4][6] <= 18'd0;\
                conv1_result[5][4][7] <= 18'd0;\
                conv1_result[5][4][8] <= 18'd0;\
                conv1_result[5][4][9] <= 18'd0;\
                conv1_result[5][4][10] <= 18'd0;\
                conv1_result[5][4][11] <= 18'd0;\
                conv1_result[5][4][12] <= 18'd0;\
                conv1_result[5][4][13] <= 18'd0;\
                conv1_result[5][5][0] <= 18'd0;\
                conv1_result[5][5][1] <= 18'd0;\
                conv1_result[5][5][2] <= 18'd0;\
                conv1_result[5][5][3] <= 18'd0;\
                conv1_result[5][5][4] <= 18'd0;\
                conv1_result[5][5][5] <= 18'd0;\
                conv1_result[5][5][6] <= 18'd0;\
                conv1_result[5][5][7] <= 18'd0;\
                conv1_result[5][5][8] <= 18'd0;\
                conv1_result[5][5][9] <= 18'd0;\
                conv1_result[5][5][10] <= 18'd0;\
                conv1_result[5][5][11] <= 18'd0;\
                conv1_result[5][5][12] <= 18'd0;\
                conv1_result[5][5][13] <= 18'd0;\
                conv1_result[5][6][0] <= 18'd0;\
                conv1_result[5][6][1] <= 18'd0;\
                conv1_result[5][6][2] <= 18'd0;\
                conv1_result[5][6][3] <= 18'd0;\
                conv1_result[5][6][4] <= 18'd0;\
                conv1_result[5][6][5] <= 18'd0;\
                conv1_result[5][6][6] <= 18'd0;\
                conv1_result[5][6][7] <= 18'd0;\
                conv1_result[5][6][8] <= 18'd0;\
                conv1_result[5][6][9] <= 18'd0;\
                conv1_result[5][6][10] <= 18'd0;\
                conv1_result[5][6][11] <= 18'd0;\
                conv1_result[5][6][12] <= 18'd0;\
                conv1_result[5][6][13] <= 18'd0;\
                conv1_result[5][7][0] <= 18'd0;\
                conv1_result[5][7][1] <= 18'd0;\
                conv1_result[5][7][2] <= 18'd0;\
                conv1_result[5][7][3] <= 18'd0;\
                conv1_result[5][7][4] <= 18'd0;\
                conv1_result[5][7][5] <= 18'd0;\
                conv1_result[5][7][6] <= 18'd0;\
                conv1_result[5][7][7] <= 18'd0;\
                conv1_result[5][7][8] <= 18'd0;\
                conv1_result[5][7][9] <= 18'd0;\
                conv1_result[5][7][10] <= 18'd0;\
                conv1_result[5][7][11] <= 18'd0;\
                conv1_result[5][7][12] <= 18'd0;\
                conv1_result[5][7][13] <= 18'd0;\
                conv1_result[5][8][0] <= 18'd0;\
                conv1_result[5][8][1] <= 18'd0;\
                conv1_result[5][8][2] <= 18'd0;\
                conv1_result[5][8][3] <= 18'd0;\
                conv1_result[5][8][4] <= 18'd0;\
                conv1_result[5][8][5] <= 18'd0;\
                conv1_result[5][8][6] <= 18'd0;\
                conv1_result[5][8][7] <= 18'd0;\
                conv1_result[5][8][8] <= 18'd0;\
                conv1_result[5][8][9] <= 18'd0;\
                conv1_result[5][8][10] <= 18'd0;\
                conv1_result[5][8][11] <= 18'd0;\
                conv1_result[5][8][12] <= 18'd0;\
                conv1_result[5][8][13] <= 18'd0;\
                conv1_result[5][9][0] <= 18'd0;\
                conv1_result[5][9][1] <= 18'd0;\
                conv1_result[5][9][2] <= 18'd0;\
                conv1_result[5][9][3] <= 18'd0;\
                conv1_result[5][9][4] <= 18'd0;\
                conv1_result[5][9][5] <= 18'd0;\
                conv1_result[5][9][6] <= 18'd0;\
                conv1_result[5][9][7] <= 18'd0;\
                conv1_result[5][9][8] <= 18'd0;\
                conv1_result[5][9][9] <= 18'd0;\
                conv1_result[5][9][10] <= 18'd0;\
                conv1_result[5][9][11] <= 18'd0;\
                conv1_result[5][9][12] <= 18'd0;\
                conv1_result[5][9][13] <= 18'd0;\
                conv1_result[5][10][0] <= 18'd0;\
                conv1_result[5][10][1] <= 18'd0;\
                conv1_result[5][10][2] <= 18'd0;\
                conv1_result[5][10][3] <= 18'd0;\
                conv1_result[5][10][4] <= 18'd0;\
                conv1_result[5][10][5] <= 18'd0;\
                conv1_result[5][10][6] <= 18'd0;\
                conv1_result[5][10][7] <= 18'd0;\
                conv1_result[5][10][8] <= 18'd0;\
                conv1_result[5][10][9] <= 18'd0;\
                conv1_result[5][10][10] <= 18'd0;\
                conv1_result[5][10][11] <= 18'd0;\
                conv1_result[5][10][12] <= 18'd0;\
                conv1_result[5][10][13] <= 18'd0;\
                conv1_result[5][11][0] <= 18'd0;\
                conv1_result[5][11][1] <= 18'd0;\
                conv1_result[5][11][2] <= 18'd0;\
                conv1_result[5][11][3] <= 18'd0;\
                conv1_result[5][11][4] <= 18'd0;\
                conv1_result[5][11][5] <= 18'd0;\
                conv1_result[5][11][6] <= 18'd0;\
                conv1_result[5][11][7] <= 18'd0;\
                conv1_result[5][11][8] <= 18'd0;\
                conv1_result[5][11][9] <= 18'd0;\
                conv1_result[5][11][10] <= 18'd0;\
                conv1_result[5][11][11] <= 18'd0;\
                conv1_result[5][11][12] <= 18'd0;\
                conv1_result[5][11][13] <= 18'd0;\
                conv1_result[5][12][0] <= 18'd0;\
                conv1_result[5][12][1] <= 18'd0;\
                conv1_result[5][12][2] <= 18'd0;\
                conv1_result[5][12][3] <= 18'd0;\
                conv1_result[5][12][4] <= 18'd0;\
                conv1_result[5][12][5] <= 18'd0;\
                conv1_result[5][12][6] <= 18'd0;\
                conv1_result[5][12][7] <= 18'd0;\
                conv1_result[5][12][8] <= 18'd0;\
                conv1_result[5][12][9] <= 18'd0;\
                conv1_result[5][12][10] <= 18'd0;\
                conv1_result[5][12][11] <= 18'd0;\
                conv1_result[5][12][12] <= 18'd0;\
                conv1_result[5][12][13] <= 18'd0;\
                conv1_result[5][13][0] <= 18'd0;\
                conv1_result[5][13][1] <= 18'd0;\
                conv1_result[5][13][2] <= 18'd0;\
                conv1_result[5][13][3] <= 18'd0;\
                conv1_result[5][13][4] <= 18'd0;\
                conv1_result[5][13][5] <= 18'd0;\
                conv1_result[5][13][6] <= 18'd0;\
                conv1_result[5][13][7] <= 18'd0;\
                conv1_result[5][13][8] <= 18'd0;\
                conv1_result[5][13][9] <= 18'd0;\
                conv1_result[5][13][10] <= 18'd0;\
                conv1_result[5][13][11] <= 18'd0;\
                conv1_result[5][13][12] <= 18'd0;\
                conv1_result[5][13][13] <= 18'd0;\
            end\
            INPUT    :;\
            CONV1_1_1:;\
            CONV1_1_2:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[0][0][0] <= compare_result[0]; conv1_result[0][0][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][0][2] <= compare_result[0]; conv1_result[0][0][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][0][4] <= compare_result[0]; conv1_result[0][0][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][0][6] <= compare_result[0]; conv1_result[0][0][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][0][8] <= compare_result[0]; conv1_result[0][0][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][0][10] <= compare_result[0]; conv1_result[0][0][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][0][12] <= compare_result[0]; conv1_result[0][0][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][1][0] <= compare_result[0]; conv1_result[0][1][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][1][2] <= compare_result[0]; conv1_result[0][1][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][1][4] <= compare_result[0]; conv1_result[0][1][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][1][6] <= compare_result[0]; conv1_result[0][1][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][1][8] <= compare_result[0]; conv1_result[0][1][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][1][10] <= compare_result[0]; conv1_result[0][1][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][1][12] <= compare_result[0]; conv1_result[0][1][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_1_3:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[0][2][0] <= compare_result[0]; conv1_result[0][2][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][2][2] <= compare_result[0]; conv1_result[0][2][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][2][4] <= compare_result[0]; conv1_result[0][2][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][2][6] <= compare_result[0]; conv1_result[0][2][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][2][ 8] <= compare_result[0]; conv1_result[0][2][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][2][10] <= compare_result[0]; conv1_result[0][2][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][2][12] <= compare_result[0]; conv1_result[0][2][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][3][ 0] <= compare_result[0]; conv1_result[0][3][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][3][ 2] <= compare_result[0]; conv1_result[0][3][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][3][ 4] <= compare_result[0]; conv1_result[0][3][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][3][ 6] <= compare_result[0]; conv1_result[0][3][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][3][ 8] <= compare_result[0]; conv1_result[0][3][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][3][10] <= compare_result[0]; conv1_result[0][3][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][3][12] <= compare_result[0]; conv1_result[0][3][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_1_4:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[0][4][ 0] <= compare_result[0]; conv1_result[0][4][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][4][ 2] <= compare_result[0]; conv1_result[0][4][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][4][ 4] <= compare_result[0]; conv1_result[0][4][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][4][ 6] <= compare_result[0]; conv1_result[0][4][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][4][ 8] <= compare_result[0]; conv1_result[0][4][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][4][10] <= compare_result[0]; conv1_result[0][4][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][4][12] <= compare_result[0]; conv1_result[0][4][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][5][ 0] <= compare_result[0]; conv1_result[0][5][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][5][ 2] <= compare_result[0]; conv1_result[0][5][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][5][ 4] <= compare_result[0]; conv1_result[0][5][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][5][ 6] <= compare_result[0]; conv1_result[0][5][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][5][ 8] <= compare_result[0]; conv1_result[0][5][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][5][10] <= compare_result[0]; conv1_result[0][5][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][5][12] <= compare_result[0]; conv1_result[0][5][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_1_5:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[0][6][ 0] <= compare_result[0]; conv1_result[0][6][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][6][ 2] <= compare_result[0]; conv1_result[0][6][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][6][ 4] <= compare_result[0]; conv1_result[0][6][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][6][ 6] <= compare_result[0]; conv1_result[0][6][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][6][ 8] <= compare_result[0]; conv1_result[0][6][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][6][10] <= compare_result[0]; conv1_result[0][6][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][6][12] <= compare_result[0]; conv1_result[0][6][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][7][ 0] <= compare_result[0]; conv1_result[0][7][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][7][ 2] <= compare_result[0]; conv1_result[0][7][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][7][ 4] <= compare_result[0]; conv1_result[0][7][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][7][ 6] <= compare_result[0]; conv1_result[0][7][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][7][ 8] <= compare_result[0]; conv1_result[0][7][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][7][10] <= compare_result[0]; conv1_result[0][7][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][7][12] <= compare_result[0]; conv1_result[0][7][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_1_6:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[0][8][ 0] <= compare_result[0]; conv1_result[0][8][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][8][ 2] <= compare_result[0]; conv1_result[0][8][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][8][ 4] <= compare_result[0]; conv1_result[0][8][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][8][ 6] <= compare_result[0]; conv1_result[0][8][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][8][ 8] <= compare_result[0]; conv1_result[0][8][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][8][10] <= compare_result[0]; conv1_result[0][8][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][8][12] <= compare_result[0]; conv1_result[0][8][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][9][ 0] <= compare_result[0]; conv1_result[0][9][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][9][ 2] <= compare_result[0]; conv1_result[0][9][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][9][ 4] <= compare_result[0]; conv1_result[0][9][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][9][ 6] <= compare_result[0]; conv1_result[0][9][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][9][ 8] <= compare_result[0]; conv1_result[0][9][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][9][10] <= compare_result[0]; conv1_result[0][9][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][9][12] <= compare_result[0]; conv1_result[0][9][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_1_7:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[0][10][ 0] <= compare_result[0]; conv1_result[0][10][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][10][ 2] <= compare_result[0]; conv1_result[0][10][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][10][ 4] <= compare_result[0]; conv1_result[0][10][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][10][ 6] <= compare_result[0]; conv1_result[0][10][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][10][ 8] <= compare_result[0]; conv1_result[0][10][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][10][10] <= compare_result[0]; conv1_result[0][10][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][10][12] <= compare_result[0]; conv1_result[0][10][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][11][ 0] <= compare_result[0]; conv1_result[0][11][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][11][ 2] <= compare_result[0]; conv1_result[0][11][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][11][ 4] <= compare_result[0]; conv1_result[0][11][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][11][ 6] <= compare_result[0]; conv1_result[0][11][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][11][ 8] <= compare_result[0]; conv1_result[0][11][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][11][10] <= compare_result[0]; conv1_result[0][11][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][11][12] <= compare_result[0]; conv1_result[0][11][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_2_1:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[0][12][ 0] <= compare_result[0]; conv1_result[0][12][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][12][ 2] <= compare_result[0]; conv1_result[0][12][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][12][ 4] <= compare_result[0]; conv1_result[0][12][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][12][ 6] <= compare_result[0]; conv1_result[0][12][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][12][ 8] <= compare_result[0]; conv1_result[0][12][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][12][10] <= compare_result[0]; conv1_result[0][12][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][12][12] <= compare_result[0]; conv1_result[0][12][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][13][ 0] <= compare_result[0]; conv1_result[0][13][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][13][ 2] <= compare_result[0]; conv1_result[0][13][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[0][13][ 4] <= compare_result[0]; conv1_result[0][13][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[0][13][ 6] <= compare_result[0]; conv1_result[0][13][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[0][13][ 8] <= compare_result[0]; conv1_result[0][13][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[0][13][10] <= compare_result[0]; conv1_result[0][13][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[0][13][12] <= compare_result[0]; conv1_result[0][13][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_2_2:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[1][ 0][ 0] <= compare_result[0]; conv1_result[1][0][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 0][ 2] <= compare_result[0]; conv1_result[1][0][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 0][ 4] <= compare_result[0]; conv1_result[1][0][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 0][ 6] <= compare_result[0]; conv1_result[1][0][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 0][ 8] <= compare_result[0]; conv1_result[1][0][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 0][10] <= compare_result[0]; conv1_result[1][0][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 0][12] <= compare_result[0]; conv1_result[1][0][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 1][ 0] <= compare_result[0]; conv1_result[1][1][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 1][ 2] <= compare_result[0]; conv1_result[1][1][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 1][ 4] <= compare_result[0]; conv1_result[1][1][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 1][ 6] <= compare_result[0]; conv1_result[1][1][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 1][ 8] <= compare_result[0]; conv1_result[1][1][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 1][10] <= compare_result[0]; conv1_result[1][1][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 1][12] <= compare_result[0]; conv1_result[1][1][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_2_3:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[1][ 2][ 0] <= compare_result[0]; conv1_result[1][2][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 2][ 2] <= compare_result[0]; conv1_result[1][2][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 2][ 4] <= compare_result[0]; conv1_result[1][2][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 2][ 6] <= compare_result[0]; conv1_result[1][2][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 2][ 8] <= compare_result[0]; conv1_result[1][2][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 2][10] <= compare_result[0]; conv1_result[1][2][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 2][12] <= compare_result[0]; conv1_result[1][2][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 3][ 0] <= compare_result[0]; conv1_result[1][3][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 3][ 2] <= compare_result[0]; conv1_result[1][3][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 3][ 4] <= compare_result[0]; conv1_result[1][3][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 3][ 6] <= compare_result[0]; conv1_result[1][3][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 3][ 8] <= compare_result[0]; conv1_result[1][3][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 3][10] <= compare_result[0]; conv1_result[1][3][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 3][12] <= compare_result[0]; conv1_result[1][3][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_2_4:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[1][ 4][ 0] <= compare_result[0]; conv1_result[1][4][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 4][ 2] <= compare_result[0]; conv1_result[1][4][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 4][ 4] <= compare_result[0]; conv1_result[1][4][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 4][ 6] <= compare_result[0]; conv1_result[1][4][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 4][ 8] <= compare_result[0]; conv1_result[1][4][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 4][10] <= compare_result[0]; conv1_result[1][4][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 4][12] <= compare_result[0]; conv1_result[1][4][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 5][ 0] <= compare_result[0]; conv1_result[1][5][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 5][ 2] <= compare_result[0]; conv1_result[1][5][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 5][ 4] <= compare_result[0]; conv1_result[1][5][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 5][ 6] <= compare_result[0]; conv1_result[1][5][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 5][ 8] <= compare_result[0]; conv1_result[1][5][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 5][10] <= compare_result[0]; conv1_result[1][5][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 5][12] <= compare_result[0]; conv1_result[1][5][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_2_5:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[1][ 6][ 0] <= compare_result[0]; conv1_result[1][6][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 6][ 2] <= compare_result[0]; conv1_result[1][6][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 6][ 4] <= compare_result[0]; conv1_result[1][6][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 6][ 6] <= compare_result[0]; conv1_result[1][6][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 6][ 8] <= compare_result[0]; conv1_result[1][6][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 6][10] <= compare_result[0]; conv1_result[1][6][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 6][12] <= compare_result[0]; conv1_result[1][6][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 7][ 0] <= compare_result[0]; conv1_result[1][7][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 7][ 2] <= compare_result[0]; conv1_result[1][7][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 7][ 4] <= compare_result[0]; conv1_result[1][7][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 7][ 6] <= compare_result[0]; conv1_result[1][7][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 7][ 8] <= compare_result[0]; conv1_result[1][7][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 7][10] <= compare_result[0]; conv1_result[1][7][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 7][12] <= compare_result[0]; conv1_result[1][7][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_2_6:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[1][ 8][ 0] <= compare_result[0]; conv1_result[1][8][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 8][ 2] <= compare_result[0]; conv1_result[1][8][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 8][ 4] <= compare_result[0]; conv1_result[1][8][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 8][ 6] <= compare_result[0]; conv1_result[1][8][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 8][ 8] <= compare_result[0]; conv1_result[1][8][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 8][10] <= compare_result[0]; conv1_result[1][8][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 8][12] <= compare_result[0]; conv1_result[1][8][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 9][ 0] <= compare_result[0]; conv1_result[1][9][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 9][ 2] <= compare_result[0]; conv1_result[1][9][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][ 9][ 4] <= compare_result[0]; conv1_result[1][9][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][ 9][ 6] <= compare_result[0]; conv1_result[1][9][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][ 9][ 8] <= compare_result[0]; conv1_result[1][9][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][ 9][10] <= compare_result[0]; conv1_result[1][9][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][ 9][12] <= compare_result[0]; conv1_result[1][9][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_2_7:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[1][10][ 0] <= compare_result[0]; conv1_result[1][10][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][10][ 2] <= compare_result[0]; conv1_result[1][10][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][10][ 4] <= compare_result[0]; conv1_result[1][10][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][10][ 6] <= compare_result[0]; conv1_result[1][10][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][10][ 8] <= compare_result[0]; conv1_result[1][10][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][10][10] <= compare_result[0]; conv1_result[1][10][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][10][12] <= compare_result[0]; conv1_result[1][10][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][11][ 0] <= compare_result[0]; conv1_result[1][11][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][11][ 2] <= compare_result[0]; conv1_result[1][11][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][11][ 4] <= compare_result[0]; conv1_result[1][11][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][11][ 6] <= compare_result[0]; conv1_result[1][11][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][11][ 8] <= compare_result[0]; conv1_result[1][11][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][11][10] <= compare_result[0]; conv1_result[1][11][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][11][12] <= compare_result[0]; conv1_result[1][11][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_3_1:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[1][12][ 0] <= compare_result[0]; conv1_result[1][12][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][12][ 2] <= compare_result[0]; conv1_result[1][12][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][12][ 4] <= compare_result[0]; conv1_result[1][12][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][12][ 6] <= compare_result[0]; conv1_result[1][12][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][12][ 8] <= compare_result[0]; conv1_result[1][12][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][12][10] <= compare_result[0]; conv1_result[1][12][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][12][12] <= compare_result[0]; conv1_result[1][12][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][13][ 0] <= compare_result[0]; conv1_result[1][13][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][13][ 2] <= compare_result[0]; conv1_result[1][13][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[1][13][ 4] <= compare_result[0]; conv1_result[1][13][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[1][13][ 6] <= compare_result[0]; conv1_result[1][13][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[1][13][ 8] <= compare_result[0]; conv1_result[1][13][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[1][13][10] <= compare_result[0]; conv1_result[1][13][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[1][13][12] <= compare_result[0]; conv1_result[1][13][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_3_2:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[2][ 0][ 0] <= compare_result[0]; conv1_result[2][0][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 0][ 2] <= compare_result[0]; conv1_result[2][0][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 0][ 4] <= compare_result[0]; conv1_result[2][0][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 0][ 6] <= compare_result[0]; conv1_result[2][0][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 0][ 8] <= compare_result[0]; conv1_result[2][0][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 0][10] <= compare_result[0]; conv1_result[2][0][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 0][12] <= compare_result[0]; conv1_result[2][0][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 1][ 0] <= compare_result[0]; conv1_result[2][1][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 1][ 2] <= compare_result[0]; conv1_result[2][1][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 1][ 4] <= compare_result[0]; conv1_result[2][1][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 1][ 6] <= compare_result[0]; conv1_result[2][1][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 1][ 8] <= compare_result[0]; conv1_result[2][1][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 1][10] <= compare_result[0]; conv1_result[2][1][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 1][12] <= compare_result[0]; conv1_result[2][1][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_3_3:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[2][ 2][ 0] <= compare_result[0]; conv1_result[2][2][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 2][ 2] <= compare_result[0]; conv1_result[2][2][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 2][ 4] <= compare_result[0]; conv1_result[2][2][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 2][ 6] <= compare_result[0]; conv1_result[2][2][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 2][ 8] <= compare_result[0]; conv1_result[2][2][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 2][10] <= compare_result[0]; conv1_result[2][2][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 2][12] <= compare_result[0]; conv1_result[2][2][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 3][ 0] <= compare_result[0]; conv1_result[2][3][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 3][ 2] <= compare_result[0]; conv1_result[2][3][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 3][ 4] <= compare_result[0]; conv1_result[2][3][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 3][ 6] <= compare_result[0]; conv1_result[2][3][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 3][ 8] <= compare_result[0]; conv1_result[2][3][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 3][10] <= compare_result[0]; conv1_result[2][3][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 3][12] <= compare_result[0]; conv1_result[2][3][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_3_4:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[2][ 4][ 0] <= compare_result[0]; conv1_result[2][4][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 4][ 2] <= compare_result[0]; conv1_result[2][4][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 4][ 4] <= compare_result[0]; conv1_result[2][4][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 4][ 6] <= compare_result[0]; conv1_result[2][4][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 4][ 8] <= compare_result[0]; conv1_result[2][4][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 4][10] <= compare_result[0]; conv1_result[2][4][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 4][12] <= compare_result[0]; conv1_result[2][4][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 5][ 0] <= compare_result[0]; conv1_result[2][5][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 5][ 2] <= compare_result[0]; conv1_result[2][5][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 5][ 4] <= compare_result[0]; conv1_result[2][5][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 5][ 6] <= compare_result[0]; conv1_result[2][5][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 5][ 8] <= compare_result[0]; conv1_result[2][5][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 5][10] <= compare_result[0]; conv1_result[2][5][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 5][12] <= compare_result[0]; conv1_result[2][5][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_3_5:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[2][ 6][ 0] <= compare_result[0]; conv1_result[2][6][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 6][ 2] <= compare_result[0]; conv1_result[2][6][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 6][ 4] <= compare_result[0]; conv1_result[2][6][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 6][ 6] <= compare_result[0]; conv1_result[2][6][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 6][ 8] <= compare_result[0]; conv1_result[2][6][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 6][10] <= compare_result[0]; conv1_result[2][6][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 6][12] <= compare_result[0]; conv1_result[2][6][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 7][ 0] <= compare_result[0]; conv1_result[2][7][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 7][ 2] <= compare_result[0]; conv1_result[2][7][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 7][ 4] <= compare_result[0]; conv1_result[2][7][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 7][ 6] <= compare_result[0]; conv1_result[2][7][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 7][ 8] <= compare_result[0]; conv1_result[2][7][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 7][10] <= compare_result[0]; conv1_result[2][7][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 7][12] <= compare_result[0]; conv1_result[2][7][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_3_6:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[2][ 8][ 0] <= compare_result[0]; conv1_result[2][8][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 8][ 2] <= compare_result[0]; conv1_result[2][8][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 8][ 4] <= compare_result[0]; conv1_result[2][8][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 8][ 6] <= compare_result[0]; conv1_result[2][8][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 8][ 8] <= compare_result[0]; conv1_result[2][8][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 8][10] <= compare_result[0]; conv1_result[2][8][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 8][12] <= compare_result[0]; conv1_result[2][8][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 9][ 0] <= compare_result[0]; conv1_result[2][9][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 9][ 2] <= compare_result[0]; conv1_result[2][9][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][ 9][ 4] <= compare_result[0]; conv1_result[2][9][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][ 9][ 6] <= compare_result[0]; conv1_result[2][9][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][ 9][ 8] <= compare_result[0]; conv1_result[2][9][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][ 9][10] <= compare_result[0]; conv1_result[2][9][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][ 9][12] <= compare_result[0]; conv1_result[2][9][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_3_7:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[2][10][ 0] <= compare_result[0]; conv1_result[2][10][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][10][ 2] <= compare_result[0]; conv1_result[2][10][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][10][ 4] <= compare_result[0]; conv1_result[2][10][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][10][ 6] <= compare_result[0]; conv1_result[2][10][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][10][ 8] <= compare_result[0]; conv1_result[2][10][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][10][10] <= compare_result[0]; conv1_result[2][10][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][10][12] <= compare_result[0]; conv1_result[2][10][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][11][ 0] <= compare_result[0]; conv1_result[2][11][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][11][ 2] <= compare_result[0]; conv1_result[2][11][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][11][ 4] <= compare_result[0]; conv1_result[2][11][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][11][ 6] <= compare_result[0]; conv1_result[2][11][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][11][ 8] <= compare_result[0]; conv1_result[2][11][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][11][10] <= compare_result[0]; conv1_result[2][11][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][11][12] <= compare_result[0]; conv1_result[2][11][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_4_1:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[2][12][ 0] <= compare_result[0]; conv1_result[2][12][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][12][ 2] <= compare_result[0]; conv1_result[2][12][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][12][ 4] <= compare_result[0]; conv1_result[2][12][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][12][ 6] <= compare_result[0]; conv1_result[2][12][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][12][ 8] <= compare_result[0]; conv1_result[2][12][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][12][10] <= compare_result[0]; conv1_result[2][12][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][12][12] <= compare_result[0]; conv1_result[2][12][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][13][ 0] <= compare_result[0]; conv1_result[2][13][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][13][ 2] <= compare_result[0]; conv1_result[2][13][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[2][13][ 4] <= compare_result[0]; conv1_result[2][13][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[2][13][ 6] <= compare_result[0]; conv1_result[2][13][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[2][13][ 8] <= compare_result[0]; conv1_result[2][13][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[2][13][10] <= compare_result[0]; conv1_result[2][13][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[2][13][12] <= compare_result[0]; conv1_result[2][13][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_4_2:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[3][ 0][ 0] <= compare_result[0]; conv1_result[3][0][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 0][ 2] <= compare_result[0]; conv1_result[3][0][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 0][ 4] <= compare_result[0]; conv1_result[3][0][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 0][ 6] <= compare_result[0]; conv1_result[3][0][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 0][ 8] <= compare_result[0]; conv1_result[3][0][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 0][10] <= compare_result[0]; conv1_result[3][0][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 0][12] <= compare_result[0]; conv1_result[3][0][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 1][ 0] <= compare_result[0]; conv1_result[3][1][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 1][ 2] <= compare_result[0]; conv1_result[3][1][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 1][ 4] <= compare_result[0]; conv1_result[3][1][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 1][ 6] <= compare_result[0]; conv1_result[3][1][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 1][ 8] <= compare_result[0]; conv1_result[3][1][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 1][10] <= compare_result[0]; conv1_result[3][1][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 1][12] <= compare_result[0]; conv1_result[3][1][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_4_3:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[3][ 2][ 0] <= compare_result[0]; conv1_result[3][2][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 2][ 2] <= compare_result[0]; conv1_result[3][2][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 2][ 4] <= compare_result[0]; conv1_result[3][2][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 2][ 6] <= compare_result[0]; conv1_result[3][2][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 2][ 8] <= compare_result[0]; conv1_result[3][2][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 2][10] <= compare_result[0]; conv1_result[3][2][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 2][12] <= compare_result[0]; conv1_result[3][2][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 3][ 0] <= compare_result[0]; conv1_result[3][3][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 3][ 2] <= compare_result[0]; conv1_result[3][3][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 3][ 4] <= compare_result[0]; conv1_result[3][3][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 3][ 6] <= compare_result[0]; conv1_result[3][3][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 3][ 8] <= compare_result[0]; conv1_result[3][3][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 3][10] <= compare_result[0]; conv1_result[3][3][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 3][12] <= compare_result[0]; conv1_result[3][3][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_4_4:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[3][ 4][ 0] <= compare_result[0]; conv1_result[3][4][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 4][ 2] <= compare_result[0]; conv1_result[3][4][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 4][ 4] <= compare_result[0]; conv1_result[3][4][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 4][ 6] <= compare_result[0]; conv1_result[3][4][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 4][ 8] <= compare_result[0]; conv1_result[3][4][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 4][10] <= compare_result[0]; conv1_result[3][4][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 4][12] <= compare_result[0]; conv1_result[3][4][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 5][ 0] <= compare_result[0]; conv1_result[3][5][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 5][ 2] <= compare_result[0]; conv1_result[3][5][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 5][ 4] <= compare_result[0]; conv1_result[3][5][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 5][ 6] <= compare_result[0]; conv1_result[3][5][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 5][ 8] <= compare_result[0]; conv1_result[3][5][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 5][10] <= compare_result[0]; conv1_result[3][5][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 5][12] <= compare_result[0]; conv1_result[3][5][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_4_5:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[3][ 6][ 0] <= compare_result[0]; conv1_result[3][6][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 6][ 2] <= compare_result[0]; conv1_result[3][6][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 6][ 4] <= compare_result[0]; conv1_result[3][6][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 6][ 6] <= compare_result[0]; conv1_result[3][6][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 6][ 8] <= compare_result[0]; conv1_result[3][6][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 6][10] <= compare_result[0]; conv1_result[3][6][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 6][12] <= compare_result[0]; conv1_result[3][6][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 7][ 0] <= compare_result[0]; conv1_result[3][7][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 7][ 2] <= compare_result[0]; conv1_result[3][7][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 7][ 4] <= compare_result[0]; conv1_result[3][7][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 7][ 6] <= compare_result[0]; conv1_result[3][7][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 7][ 8] <= compare_result[0]; conv1_result[3][7][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 7][10] <= compare_result[0]; conv1_result[3][7][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 7][12] <= compare_result[0]; conv1_result[3][7][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_4_6:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[3][ 8][ 0] <= compare_result[0]; conv1_result[3][8][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 8][ 2] <= compare_result[0]; conv1_result[3][8][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 8][ 4] <= compare_result[0]; conv1_result[3][8][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 8][ 6] <= compare_result[0]; conv1_result[3][8][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 8][ 8] <= compare_result[0]; conv1_result[3][8][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 8][10] <= compare_result[0]; conv1_result[3][8][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 8][12] <= compare_result[0]; conv1_result[3][8][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 9][ 0] <= compare_result[0]; conv1_result[3][9][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 9][ 2] <= compare_result[0]; conv1_result[3][9][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][ 9][ 4] <= compare_result[0]; conv1_result[3][9][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][ 9][ 6] <= compare_result[0]; conv1_result[3][9][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][ 9][ 8] <= compare_result[0]; conv1_result[3][9][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][ 9][10] <= compare_result[0]; conv1_result[3][9][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][ 9][12] <= compare_result[0]; conv1_result[3][9][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_4_7:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[3][10][ 0] <= compare_result[0]; conv1_result[3][10][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][10][ 2] <= compare_result[0]; conv1_result[3][10][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][10][ 4] <= compare_result[0]; conv1_result[3][10][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][10][ 6] <= compare_result[0]; conv1_result[3][10][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][10][ 8] <= compare_result[0]; conv1_result[3][10][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][10][10] <= compare_result[0]; conv1_result[3][10][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][10][12] <= compare_result[0]; conv1_result[3][10][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][11][ 0] <= compare_result[0]; conv1_result[3][11][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][11][ 2] <= compare_result[0]; conv1_result[3][11][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][11][ 4] <= compare_result[0]; conv1_result[3][11][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][11][ 6] <= compare_result[0]; conv1_result[3][11][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][11][ 8] <= compare_result[0]; conv1_result[3][11][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][11][10] <= compare_result[0]; conv1_result[3][11][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][11][12] <= compare_result[0]; conv1_result[3][11][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_5_1:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[3][12][ 0] <= compare_result[0]; conv1_result[3][12][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][12][ 2] <= compare_result[0]; conv1_result[3][12][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][12][ 4] <= compare_result[0]; conv1_result[3][12][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][12][ 6] <= compare_result[0]; conv1_result[3][12][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][12][ 8] <= compare_result[0]; conv1_result[3][12][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][12][10] <= compare_result[0]; conv1_result[3][12][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][12][12] <= compare_result[0]; conv1_result[3][12][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][13][ 0] <= compare_result[0]; conv1_result[3][13][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][13][ 2] <= compare_result[0]; conv1_result[3][13][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[3][13][ 4] <= compare_result[0]; conv1_result[3][13][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[3][13][ 6] <= compare_result[0]; conv1_result[3][13][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[3][13][ 8] <= compare_result[0]; conv1_result[3][13][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[3][13][10] <= compare_result[0]; conv1_result[3][13][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[3][13][12] <= compare_result[0]; conv1_result[3][13][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_5_2:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[4][ 0][ 0] <= compare_result[0]; conv1_result[4][0][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 0][ 2] <= compare_result[0]; conv1_result[4][0][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 0][ 4] <= compare_result[0]; conv1_result[4][0][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 0][ 6] <= compare_result[0]; conv1_result[4][0][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 0][ 8] <= compare_result[0]; conv1_result[4][0][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 0][10] <= compare_result[0]; conv1_result[4][0][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 0][12] <= compare_result[0]; conv1_result[4][0][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 1][ 0] <= compare_result[0]; conv1_result[4][1][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 1][ 2] <= compare_result[0]; conv1_result[4][1][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 1][ 4] <= compare_result[0]; conv1_result[4][1][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 1][ 6] <= compare_result[0]; conv1_result[4][1][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 1][ 8] <= compare_result[0]; conv1_result[4][1][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 1][10] <= compare_result[0]; conv1_result[4][1][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 1][12] <= compare_result[0]; conv1_result[4][1][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_5_3:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[4][ 2][ 0] <= compare_result[0]; conv1_result[4][2][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 2][ 2] <= compare_result[0]; conv1_result[4][2][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 2][ 4] <= compare_result[0]; conv1_result[4][2][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 2][ 6] <= compare_result[0]; conv1_result[4][2][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 2][ 8] <= compare_result[0]; conv1_result[4][2][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 2][10] <= compare_result[0]; conv1_result[4][2][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 2][12] <= compare_result[0]; conv1_result[4][2][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 3][ 0] <= compare_result[0]; conv1_result[4][3][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 3][ 2] <= compare_result[0]; conv1_result[4][3][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 3][ 4] <= compare_result[0]; conv1_result[4][3][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 3][ 6] <= compare_result[0]; conv1_result[4][3][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 3][ 8] <= compare_result[0]; conv1_result[4][3][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 3][10] <= compare_result[0]; conv1_result[4][3][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 3][12] <= compare_result[0]; conv1_result[4][3][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_5_4:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[4][ 4][ 0] <= compare_result[0]; conv1_result[4][4][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 4][ 2] <= compare_result[0]; conv1_result[4][4][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 4][ 4] <= compare_result[0]; conv1_result[4][4][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 4][ 6] <= compare_result[0]; conv1_result[4][4][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 4][ 8] <= compare_result[0]; conv1_result[4][4][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 4][10] <= compare_result[0]; conv1_result[4][4][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 4][12] <= compare_result[0]; conv1_result[4][4][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 5][ 0] <= compare_result[0]; conv1_result[4][5][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 5][ 2] <= compare_result[0]; conv1_result[4][5][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 5][ 4] <= compare_result[0]; conv1_result[4][5][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 5][ 6] <= compare_result[0]; conv1_result[4][5][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 5][ 8] <= compare_result[0]; conv1_result[4][5][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 5][10] <= compare_result[0]; conv1_result[4][5][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 5][12] <= compare_result[0]; conv1_result[4][5][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_5_5:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[4][ 6][ 0] <= compare_result[0]; conv1_result[4][6][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 6][ 2] <= compare_result[0]; conv1_result[4][6][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 6][ 4] <= compare_result[0]; conv1_result[4][6][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 6][ 6] <= compare_result[0]; conv1_result[4][6][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 6][ 8] <= compare_result[0]; conv1_result[4][6][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 6][10] <= compare_result[0]; conv1_result[4][6][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 6][12] <= compare_result[0]; conv1_result[4][6][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 7][ 0] <= compare_result[0]; conv1_result[4][7][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 7][ 2] <= compare_result[0]; conv1_result[4][7][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 7][ 4] <= compare_result[0]; conv1_result[4][7][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 7][ 6] <= compare_result[0]; conv1_result[4][7][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 7][ 8] <= compare_result[0]; conv1_result[4][7][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 7][10] <= compare_result[0]; conv1_result[4][7][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 7][12] <= compare_result[0]; conv1_result[4][7][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_5_6:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[4][ 8][ 0] <= compare_result[0]; conv1_result[4][8][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 8][ 2] <= compare_result[0]; conv1_result[4][8][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 8][ 4] <= compare_result[0]; conv1_result[4][8][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 8][ 6] <= compare_result[0]; conv1_result[4][8][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 8][ 8] <= compare_result[0]; conv1_result[4][8][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 8][10] <= compare_result[0]; conv1_result[4][8][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 8][12] <= compare_result[0]; conv1_result[4][8][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 9][ 0] <= compare_result[0]; conv1_result[4][9][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 9][ 2] <= compare_result[0]; conv1_result[4][9][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][ 9][ 4] <= compare_result[0]; conv1_result[4][9][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][ 9][ 6] <= compare_result[0]; conv1_result[4][9][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][ 9][ 8] <= compare_result[0]; conv1_result[4][9][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][ 9][10] <= compare_result[0]; conv1_result[4][9][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][ 9][12] <= compare_result[0]; conv1_result[4][9][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_5_7:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[4][10][ 0] <= compare_result[0]; conv1_result[4][10][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][10][ 2] <= compare_result[0]; conv1_result[4][10][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][10][ 4] <= compare_result[0]; conv1_result[4][10][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][10][ 6] <= compare_result[0]; conv1_result[4][10][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][10][ 8] <= compare_result[0]; conv1_result[4][10][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][10][10] <= compare_result[0]; conv1_result[4][10][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][10][12] <= compare_result[0]; conv1_result[4][10][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][11][ 0] <= compare_result[0]; conv1_result[4][11][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][11][ 2] <= compare_result[0]; conv1_result[4][11][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][11][ 4] <= compare_result[0]; conv1_result[4][11][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][11][ 6] <= compare_result[0]; conv1_result[4][11][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][11][ 8] <= compare_result[0]; conv1_result[4][11][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][11][10] <= compare_result[0]; conv1_result[4][11][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][11][12] <= compare_result[0]; conv1_result[4][11][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_6_1:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[4][12][ 0] <= compare_result[0]; conv1_result[4][12][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][12][ 2] <= compare_result[0]; conv1_result[4][12][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][12][ 4] <= compare_result[0]; conv1_result[4][12][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][12][ 6] <= compare_result[0]; conv1_result[4][12][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][12][ 8] <= compare_result[0]; conv1_result[4][12][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][12][10] <= compare_result[0]; conv1_result[4][12][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][12][12] <= compare_result[0]; conv1_result[4][12][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][13][ 0] <= compare_result[0]; conv1_result[4][13][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][13][ 2] <= compare_result[0]; conv1_result[4][13][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[4][13][ 4] <= compare_result[0]; conv1_result[4][13][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[4][13][ 6] <= compare_result[0]; conv1_result[4][13][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[4][13][ 8] <= compare_result[0]; conv1_result[4][13][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[4][13][10] <= compare_result[0]; conv1_result[4][13][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[4][13][12] <= compare_result[0]; conv1_result[4][13][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_6_2:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[5][ 0][ 0] <= compare_result[0]; conv1_result[5][0][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 0][ 2] <= compare_result[0]; conv1_result[5][0][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 0][ 4] <= compare_result[0]; conv1_result[5][0][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 0][ 6] <= compare_result[0]; conv1_result[5][0][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 0][ 8] <= compare_result[0]; conv1_result[5][0][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 0][10] <= compare_result[0]; conv1_result[5][0][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 0][12] <= compare_result[0]; conv1_result[5][0][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 1][ 0] <= compare_result[0]; conv1_result[5][1][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 1][ 2] <= compare_result[0]; conv1_result[5][1][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 1][ 4] <= compare_result[0]; conv1_result[5][1][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 1][ 6] <= compare_result[0]; conv1_result[5][1][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 1][ 8] <= compare_result[0]; conv1_result[5][1][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 1][10] <= compare_result[0]; conv1_result[5][1][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 1][12] <= compare_result[0]; conv1_result[5][1][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_6_3:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[5][ 2][ 0] <= compare_result[0]; conv1_result[5][2][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 2][ 2] <= compare_result[0]; conv1_result[5][2][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 2][ 4] <= compare_result[0]; conv1_result[5][2][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 2][ 6] <= compare_result[0]; conv1_result[5][2][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 2][ 8] <= compare_result[0]; conv1_result[5][2][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 2][10] <= compare_result[0]; conv1_result[5][2][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 2][12] <= compare_result[0]; conv1_result[5][2][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 3][ 0] <= compare_result[0]; conv1_result[5][3][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 3][ 2] <= compare_result[0]; conv1_result[5][3][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 3][ 4] <= compare_result[0]; conv1_result[5][3][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 3][ 6] <= compare_result[0]; conv1_result[5][3][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 3][ 8] <= compare_result[0]; conv1_result[5][3][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 3][10] <= compare_result[0]; conv1_result[5][3][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 3][12] <= compare_result[0]; conv1_result[5][3][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_6_4:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[5][ 4][ 0] <= compare_result[0]; conv1_result[5][4][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 4][ 2] <= compare_result[0]; conv1_result[5][4][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 4][ 4] <= compare_result[0]; conv1_result[5][4][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 4][ 6] <= compare_result[0]; conv1_result[5][4][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 4][ 8] <= compare_result[0]; conv1_result[5][4][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 4][10] <= compare_result[0]; conv1_result[5][4][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 4][12] <= compare_result[0]; conv1_result[5][4][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 5][ 0] <= compare_result[0]; conv1_result[5][5][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 5][ 2] <= compare_result[0]; conv1_result[5][5][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 5][ 4] <= compare_result[0]; conv1_result[5][5][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 5][ 6] <= compare_result[0]; conv1_result[5][5][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 5][ 8] <= compare_result[0]; conv1_result[5][5][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 5][10] <= compare_result[0]; conv1_result[5][5][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 5][12] <= compare_result[0]; conv1_result[5][5][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_6_5:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[5][ 6][ 0] <= compare_result[0]; conv1_result[5][6][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 6][ 2] <= compare_result[0]; conv1_result[5][6][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 6][ 4] <= compare_result[0]; conv1_result[5][6][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 6][ 6] <= compare_result[0]; conv1_result[5][6][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 6][ 8] <= compare_result[0]; conv1_result[5][6][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 6][10] <= compare_result[0]; conv1_result[5][6][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 6][12] <= compare_result[0]; conv1_result[5][6][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 7][ 0] <= compare_result[0]; conv1_result[5][7][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 7][ 2] <= compare_result[0]; conv1_result[5][7][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 7][ 4] <= compare_result[0]; conv1_result[5][7][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 7][ 6] <= compare_result[0]; conv1_result[5][7][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 7][ 8] <= compare_result[0]; conv1_result[5][7][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 7][10] <= compare_result[0]; conv1_result[5][7][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 7][12] <= compare_result[0]; conv1_result[5][7][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_6_6:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[5][ 8][ 0] <= compare_result[0]; conv1_result[5][8][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 8][ 2] <= compare_result[0]; conv1_result[5][8][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 8][ 4] <= compare_result[0]; conv1_result[5][8][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 8][ 6] <= compare_result[0]; conv1_result[5][8][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 8][ 8] <= compare_result[0]; conv1_result[5][8][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 8][10] <= compare_result[0]; conv1_result[5][8][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 8][12] <= compare_result[0]; conv1_result[5][8][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 9][ 0] <= compare_result[0]; conv1_result[5][9][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 9][ 2] <= compare_result[0]; conv1_result[5][9][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][ 9][ 4] <= compare_result[0]; conv1_result[5][9][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][ 9][ 6] <= compare_result[0]; conv1_result[5][9][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][ 9][ 8] <= compare_result[0]; conv1_result[5][9][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][ 9][10] <= compare_result[0]; conv1_result[5][9][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][ 9][12] <= compare_result[0]; conv1_result[5][9][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV1_6_7:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[5][10][ 0] <= compare_result[0]; conv1_result[5][10][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][10][ 2] <= compare_result[0]; conv1_result[5][10][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][10][ 4] <= compare_result[0]; conv1_result[5][10][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][10][ 6] <= compare_result[0]; conv1_result[5][10][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][10][ 8] <= compare_result[0]; conv1_result[5][10][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][10][10] <= compare_result[0]; conv1_result[5][10][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][10][12] <= compare_result[0]; conv1_result[5][10][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][11][ 0] <= compare_result[0]; conv1_result[5][11][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][11][ 2] <= compare_result[0]; conv1_result[5][11][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][11][ 4] <= compare_result[0]; conv1_result[5][11][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][11][ 6] <= compare_result[0]; conv1_result[5][11][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][11][ 8] <= compare_result[0]; conv1_result[5][11][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][11][10] <= compare_result[0]; conv1_result[5][11][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][11][12] <= compare_result[0]; conv1_result[5][11][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV2_1_1:begin\
                case(cnt1)\
                    8'd0:begin\
                        case(cnt2)\
                            8'd1:begin conv1_result[5][12][ 0] <= compare_result[0]; conv1_result[5][12][1] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][12][ 2] <= compare_result[0]; conv1_result[5][12][3] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][12][ 4] <= compare_result[0]; conv1_result[5][12][5] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][12][ 6] <= compare_result[0]; conv1_result[5][12][7] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd1:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][12][ 8] <= compare_result[0]; conv1_result[5][12][9] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][12][10] <= compare_result[0]; conv1_result[5][12][11] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][12][12] <= compare_result[0]; conv1_result[5][12][13] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][13][ 0] <= compare_result[0]; conv1_result[5][13][1] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][13][ 2] <= compare_result[0]; conv1_result[5][13][3] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    8'd2:begin\
                        case(cnt2)\
                            8'd0:begin conv1_result[5][13][ 4] <= compare_result[0]; conv1_result[5][13][5] <= compare_result[1]; end\
                            8'd1:begin conv1_result[5][13][ 6] <= compare_result[0]; conv1_result[5][13][7] <= compare_result[1]; end\
                            8'd2:begin conv1_result[5][13][ 8] <= compare_result[0]; conv1_result[5][13][9] <= compare_result[1]; end\
                            8'd3:begin conv1_result[5][13][10] <= compare_result[0]; conv1_result[5][13][11] <= compare_result[1]; end\
                            8'd4:begin conv1_result[5][13][12] <= compare_result[0]; conv1_result[5][13][13] <= compare_result[1]; end\
                            default:;\
                        endcase\
                    end\
                    default:;\
                endcase\
            end\
            CONV2_1_2,CONV2_1_3,CONV2_1_4,CONV2_1_5,CONV2_1_6,CONV2_2_1,CONV2_2_2,CONV2_2_3,CONV2_2_4,CONV2_2_5,CONV2_2_6,CONV2_3_1,CONV2_3_2,CONV2_3_3,\
            CONV2_3_4,CONV2_3_5,CONV2_3_6,CONV2_4_1,CONV2_4_2,CONV2_4_3,CONV2_4_4,CONV2_4_5,CONV2_4_6,CONV2_5_1,CONV2_5_2,CONV2_5_3,CONV2_5_4,CONV2_5_5,\
            CONV2_5_6,CONV2_6_1,CONV2_6_2,CONV2_6_3,CONV2_6_4,CONV2_6_5,CONV2_6_6,LINEAR1,LINEAR2,COMPARE,COMPLETE:;\
            default:;\
        endcase\
    end\
end