`define LINEAR1_WEIGHT \
reg [0:17] linear1_weight_array [0:11][0:149];\
always@(posedge clk) begin\
    linear1_weight_array[0][0] <= 18'h2000e;\
    linear1_weight_array[0][1] <= 18'h000cb;\
    linear1_weight_array[0][2] <= 18'h001b0;\
    linear1_weight_array[0][3] <= 18'h000d9;\
    linear1_weight_array[0][4] <= 18'h00083;\
    linear1_weight_array[0][5] <= 18'h0000d;\
    linear1_weight_array[0][6] <= 18'h001a5;\
    linear1_weight_array[0][7] <= 18'h00089;\
    linear1_weight_array[0][8] <= 18'h0004b;\
    linear1_weight_array[0][9] <= 18'h0010d;\
    linear1_weight_array[0][10] <= 18'h00095;\
    linear1_weight_array[0][11] <= 18'h000ee;\
    linear1_weight_array[0][12] <= 18'h20032;\
    linear1_weight_array[0][13] <= 18'h0013d;\
    linear1_weight_array[0][14] <= 18'h20037;\
    linear1_weight_array[0][15] <= 18'h200ad;\
    linear1_weight_array[0][16] <= 18'h20088;\
    linear1_weight_array[0][17] <= 18'h20065;\
    linear1_weight_array[0][18] <= 18'h00019;\
    linear1_weight_array[0][19] <= 18'h200c8;\
    linear1_weight_array[0][20] <= 18'h20099;\
    linear1_weight_array[0][21] <= 18'h20034;\
    linear1_weight_array[0][22] <= 18'h201b9;\
    linear1_weight_array[0][23] <= 18'h20178;\
    linear1_weight_array[0][24] <= 18'h20183;\
    linear1_weight_array[0][25] <= 18'h0007c;\
    linear1_weight_array[0][26] <= 18'h200e9;\
    linear1_weight_array[0][27] <= 18'h000ad;\
    linear1_weight_array[0][28] <= 18'h000e6;\
    linear1_weight_array[0][29] <= 18'h000e6;\
    linear1_weight_array[0][30] <= 18'h0011d;\
    linear1_weight_array[0][31] <= 18'h200a1;\
    linear1_weight_array[0][32] <= 18'h2006b;\
    linear1_weight_array[0][33] <= 18'h2005e;\
    linear1_weight_array[0][34] <= 18'h20023;\
    linear1_weight_array[0][35] <= 18'h0009b;\
    linear1_weight_array[0][36] <= 18'h0004b;\
    linear1_weight_array[0][37] <= 18'h000c0;\
    linear1_weight_array[0][38] <= 18'h2004f;\
    linear1_weight_array[0][39] <= 18'h0014d;\
    linear1_weight_array[0][40] <= 18'h00082;\
    linear1_weight_array[0][41] <= 18'h00024;\
    linear1_weight_array[0][42] <= 18'h200e8;\
    linear1_weight_array[0][43] <= 18'h20191;\
    linear1_weight_array[0][44] <= 18'h00083;\
    linear1_weight_array[0][45] <= 18'h0004b;\
    linear1_weight_array[0][46] <= 18'h20059;\
    linear1_weight_array[0][47] <= 18'h200cf;\
    linear1_weight_array[0][48] <= 18'h20030;\
    linear1_weight_array[0][49] <= 18'h000f2;\
    linear1_weight_array[0][50] <= 18'h2018f;\
    linear1_weight_array[0][51] <= 18'h2005e;\
    linear1_weight_array[0][52] <= 18'h2011d;\
    linear1_weight_array[0][53] <= 18'h200fb;\
    linear1_weight_array[0][54] <= 18'h200c0;\
    linear1_weight_array[0][55] <= 18'h2000d;\
    linear1_weight_array[0][56] <= 18'h2005b;\
    linear1_weight_array[0][57] <= 18'h0006d;\
    linear1_weight_array[0][58] <= 18'h00066;\
    linear1_weight_array[0][59] <= 18'h200a6;\
    linear1_weight_array[0][60] <= 18'h2012d;\
    linear1_weight_array[0][61] <= 18'h2011d;\
    linear1_weight_array[0][62] <= 18'h0002e;\
    linear1_weight_array[0][63] <= 18'h2001b;\
    linear1_weight_array[0][64] <= 18'h00034;\
    linear1_weight_array[0][65] <= 18'h20289;\
    linear1_weight_array[0][66] <= 18'h200e5;\
    linear1_weight_array[0][67] <= 18'h20020;\
    linear1_weight_array[0][68] <= 18'h200fe;\
    linear1_weight_array[0][69] <= 18'h00005;\
    linear1_weight_array[0][70] <= 18'h2020b;\
    linear1_weight_array[0][71] <= 18'h2021f;\
    linear1_weight_array[0][72] <= 18'h2007c;\
    linear1_weight_array[0][73] <= 18'h000c7;\
    linear1_weight_array[0][74] <= 18'h0002a;\
    linear1_weight_array[0][75] <= 18'h001c0;\
    linear1_weight_array[0][76] <= 18'h000d6;\
    linear1_weight_array[0][77] <= 18'h000a4;\
    linear1_weight_array[0][78] <= 18'h20047;\
    linear1_weight_array[0][79] <= 18'h200be;\
    linear1_weight_array[0][80] <= 18'h00077;\
    linear1_weight_array[0][81] <= 18'h2002c;\
    linear1_weight_array[0][82] <= 18'h00054;\
    linear1_weight_array[0][83] <= 18'h20042;\
    linear1_weight_array[0][84] <= 18'h20264;\
    linear1_weight_array[0][85] <= 18'h2008e;\
    linear1_weight_array[0][86] <= 18'h000c8;\
    linear1_weight_array[0][87] <= 18'h00061;\
    linear1_weight_array[0][88] <= 18'h2007f;\
    linear1_weight_array[0][89] <= 18'h20053;\
    linear1_weight_array[0][90] <= 18'h0004a;\
    linear1_weight_array[0][91] <= 18'h000ad;\
    linear1_weight_array[0][92] <= 18'h00016;\
    linear1_weight_array[0][93] <= 18'h2004c;\
    linear1_weight_array[0][94] <= 18'h200ca;\
    linear1_weight_array[0][95] <= 18'h0003a;\
    linear1_weight_array[0][96] <= 18'h0011e;\
    linear1_weight_array[0][97] <= 18'h0007a;\
    linear1_weight_array[0][98] <= 18'h001e2;\
    linear1_weight_array[0][99] <= 18'h00234;\
    linear1_weight_array[0][100] <= 18'h20193;\
    linear1_weight_array[0][101] <= 18'h2000b;\
    linear1_weight_array[0][102] <= 18'h000f3;\
    linear1_weight_array[0][103] <= 18'h0001c;\
    linear1_weight_array[0][104] <= 18'h002ea;\
    linear1_weight_array[0][105] <= 18'h000a5;\
    linear1_weight_array[0][106] <= 18'h00118;\
    linear1_weight_array[0][107] <= 18'h2006a;\
    linear1_weight_array[0][108] <= 18'h0016c;\
    linear1_weight_array[0][109] <= 18'h00095;\
    linear1_weight_array[0][110] <= 18'h0001a;\
    linear1_weight_array[0][111] <= 18'h000ac;\
    linear1_weight_array[0][112] <= 18'h00055;\
    linear1_weight_array[0][113] <= 18'h000ea;\
    linear1_weight_array[0][114] <= 18'h0008b;\
    linear1_weight_array[0][115] <= 18'h2002c;\
    linear1_weight_array[0][116] <= 18'h00107;\
    linear1_weight_array[0][117] <= 18'h001da;\
    linear1_weight_array[0][118] <= 18'h00048;\
    linear1_weight_array[0][119] <= 18'h0004c;\
    linear1_weight_array[0][120] <= 18'h2005d;\
    linear1_weight_array[0][121] <= 18'h00157;\
    linear1_weight_array[0][122] <= 18'h00118;\
    linear1_weight_array[0][123] <= 18'h2002d;\
    linear1_weight_array[0][124] <= 18'h2022d;\
    linear1_weight_array[0][125] <= 18'h000b9;\
    linear1_weight_array[0][126] <= 18'h001f4;\
    linear1_weight_array[0][127] <= 18'h00109;\
    linear1_weight_array[0][128] <= 18'h00072;\
    linear1_weight_array[0][129] <= 18'h2009e;\
    linear1_weight_array[0][130] <= 18'h000eb;\
    linear1_weight_array[0][131] <= 18'h2003a;\
    linear1_weight_array[0][132] <= 18'h0010a;\
    linear1_weight_array[0][133] <= 18'h001f9;\
    linear1_weight_array[0][134] <= 18'h20083;\
    linear1_weight_array[0][135] <= 18'h2004a;\
    linear1_weight_array[0][136] <= 18'h00098;\
    linear1_weight_array[0][137] <= 18'h000d1;\
    linear1_weight_array[0][138] <= 18'h2002c;\
    linear1_weight_array[0][139] <= 18'h20041;\
    linear1_weight_array[0][140] <= 18'h00016;\
    linear1_weight_array[0][141] <= 18'h00116;\
    linear1_weight_array[0][142] <= 18'h20053;\
    linear1_weight_array[0][143] <= 18'h20000;\
    linear1_weight_array[0][144] <= 18'h20018;\
    linear1_weight_array[0][145] <= 18'h20040;\
    linear1_weight_array[0][146] <= 18'h0010d;\
    linear1_weight_array[0][147] <= 18'h000b5;\
    linear1_weight_array[0][148] <= 18'h2007e;\
    linear1_weight_array[0][149] <= 18'h0000c;\
    linear1_weight_array[1][0] <= 18'h00004;\
    linear1_weight_array[1][1] <= 18'h0000d;\
    linear1_weight_array[1][2] <= 18'h00013;\
    linear1_weight_array[1][3] <= 18'h00011;\
    linear1_weight_array[1][4] <= 18'h2006a;\
    linear1_weight_array[1][5] <= 18'h2004d;\
    linear1_weight_array[1][6] <= 18'h0001f;\
    linear1_weight_array[1][7] <= 18'h2002b;\
    linear1_weight_array[1][8] <= 18'h0000c;\
    linear1_weight_array[1][9] <= 18'h2004b;\
    linear1_weight_array[1][10] <= 18'h00029;\
    linear1_weight_array[1][11] <= 18'h2003a;\
    linear1_weight_array[1][12] <= 18'h2002f;\
    linear1_weight_array[1][13] <= 18'h20015;\
    linear1_weight_array[1][14] <= 18'h00024;\
    linear1_weight_array[1][15] <= 18'h00019;\
    linear1_weight_array[1][16] <= 18'h00024;\
    linear1_weight_array[1][17] <= 18'h00007;\
    linear1_weight_array[1][18] <= 18'h20040;\
    linear1_weight_array[1][19] <= 18'h00036;\
    linear1_weight_array[1][20] <= 18'h20034;\
    linear1_weight_array[1][21] <= 18'h00017;\
    linear1_weight_array[1][22] <= 18'h2002c;\
    linear1_weight_array[1][23] <= 18'h0000c;\
    linear1_weight_array[1][24] <= 18'h0001e;\
    linear1_weight_array[1][25] <= 18'h20005;\
    linear1_weight_array[1][26] <= 18'h2000e;\
    linear1_weight_array[1][27] <= 18'h2002a;\
    linear1_weight_array[1][28] <= 18'h2004b;\
    linear1_weight_array[1][29] <= 18'h0001f;\
    linear1_weight_array[1][30] <= 18'h20068;\
    linear1_weight_array[1][31] <= 18'h20027;\
    linear1_weight_array[1][32] <= 18'h2004b;\
    linear1_weight_array[1][33] <= 18'h00005;\
    linear1_weight_array[1][34] <= 18'h2001f;\
    linear1_weight_array[1][35] <= 18'h2002c;\
    linear1_weight_array[1][36] <= 18'h20064;\
    linear1_weight_array[1][37] <= 18'h00028;\
    linear1_weight_array[1][38] <= 18'h2005d;\
    linear1_weight_array[1][39] <= 18'h0003b;\
    linear1_weight_array[1][40] <= 18'h0001b;\
    linear1_weight_array[1][41] <= 18'h00022;\
    linear1_weight_array[1][42] <= 18'h20064;\
    linear1_weight_array[1][43] <= 18'h20036;\
    linear1_weight_array[1][44] <= 18'h20041;\
    linear1_weight_array[1][45] <= 18'h00000;\
    linear1_weight_array[1][46] <= 18'h0000c;\
    linear1_weight_array[1][47] <= 18'h20032;\
    linear1_weight_array[1][48] <= 18'h00011;\
    linear1_weight_array[1][49] <= 18'h00031;\
    linear1_weight_array[1][50] <= 18'h00019;\
    linear1_weight_array[1][51] <= 18'h20043;\
    linear1_weight_array[1][52] <= 18'h00032;\
    linear1_weight_array[1][53] <= 18'h20051;\
    linear1_weight_array[1][54] <= 18'h00000;\
    linear1_weight_array[1][55] <= 18'h2001f;\
    linear1_weight_array[1][56] <= 18'h2003f;\
    linear1_weight_array[1][57] <= 18'h2000f;\
    linear1_weight_array[1][58] <= 18'h20046;\
    linear1_weight_array[1][59] <= 18'h2001c;\
    linear1_weight_array[1][60] <= 18'h00047;\
    linear1_weight_array[1][61] <= 18'h0002c;\
    linear1_weight_array[1][62] <= 18'h00001;\
    linear1_weight_array[1][63] <= 18'h00020;\
    linear1_weight_array[1][64] <= 18'h0001d;\
    linear1_weight_array[1][65] <= 18'h0002c;\
    linear1_weight_array[1][66] <= 18'h00027;\
    linear1_weight_array[1][67] <= 18'h20039;\
    linear1_weight_array[1][68] <= 18'h2005f;\
    linear1_weight_array[1][69] <= 18'h20058;\
    linear1_weight_array[1][70] <= 18'h20053;\
    linear1_weight_array[1][71] <= 18'h20027;\
    linear1_weight_array[1][72] <= 18'h00037;\
    linear1_weight_array[1][73] <= 18'h20010;\
    linear1_weight_array[1][74] <= 18'h00021;\
    linear1_weight_array[1][75] <= 18'h00024;\
    linear1_weight_array[1][76] <= 18'h20020;\
    linear1_weight_array[1][77] <= 18'h20055;\
    linear1_weight_array[1][78] <= 18'h20076;\
    linear1_weight_array[1][79] <= 18'h2003f;\
    linear1_weight_array[1][80] <= 18'h00019;\
    linear1_weight_array[1][81] <= 18'h2006d;\
    linear1_weight_array[1][82] <= 18'h2005d;\
    linear1_weight_array[1][83] <= 18'h20043;\
    linear1_weight_array[1][84] <= 18'h20041;\
    linear1_weight_array[1][85] <= 18'h00007;\
    linear1_weight_array[1][86] <= 18'h20069;\
    linear1_weight_array[1][87] <= 18'h00018;\
    linear1_weight_array[1][88] <= 18'h20017;\
    linear1_weight_array[1][89] <= 18'h00013;\
    linear1_weight_array[1][90] <= 18'h2002f;\
    linear1_weight_array[1][91] <= 18'h20054;\
    linear1_weight_array[1][92] <= 18'h2001b;\
    linear1_weight_array[1][93] <= 18'h20043;\
    linear1_weight_array[1][94] <= 18'h2002b;\
    linear1_weight_array[1][95] <= 18'h2002c;\
    linear1_weight_array[1][96] <= 18'h20037;\
    linear1_weight_array[1][97] <= 18'h20039;\
    linear1_weight_array[1][98] <= 18'h2002e;\
    linear1_weight_array[1][99] <= 18'h00006;\
    linear1_weight_array[1][100] <= 18'h2006c;\
    linear1_weight_array[1][101] <= 18'h20047;\
    linear1_weight_array[1][102] <= 18'h00012;\
    linear1_weight_array[1][103] <= 18'h20065;\
    linear1_weight_array[1][104] <= 18'h20054;\
    linear1_weight_array[1][105] <= 18'h00017;\
    linear1_weight_array[1][106] <= 18'h0002f;\
    linear1_weight_array[1][107] <= 18'h20017;\
    linear1_weight_array[1][108] <= 18'h20035;\
    linear1_weight_array[1][109] <= 18'h00014;\
    linear1_weight_array[1][110] <= 18'h00006;\
    linear1_weight_array[1][111] <= 18'h00002;\
    linear1_weight_array[1][112] <= 18'h20010;\
    linear1_weight_array[1][113] <= 18'h2001f;\
    linear1_weight_array[1][114] <= 18'h20022;\
    linear1_weight_array[1][115] <= 18'h2005c;\
    linear1_weight_array[1][116] <= 18'h2005d;\
    linear1_weight_array[1][117] <= 18'h2005e;\
    linear1_weight_array[1][118] <= 18'h0000e;\
    linear1_weight_array[1][119] <= 18'h2000d;\
    linear1_weight_array[1][120] <= 18'h20027;\
    linear1_weight_array[1][121] <= 18'h20004;\
    linear1_weight_array[1][122] <= 18'h20052;\
    linear1_weight_array[1][123] <= 18'h20017;\
    linear1_weight_array[1][124] <= 18'h20009;\
    linear1_weight_array[1][125] <= 18'h2001c;\
    linear1_weight_array[1][126] <= 18'h20081;\
    linear1_weight_array[1][127] <= 18'h20050;\
    linear1_weight_array[1][128] <= 18'h20044;\
    linear1_weight_array[1][129] <= 18'h00023;\
    linear1_weight_array[1][130] <= 18'h20031;\
    linear1_weight_array[1][131] <= 18'h00035;\
    linear1_weight_array[1][132] <= 18'h20057;\
    linear1_weight_array[1][133] <= 18'h2001e;\
    linear1_weight_array[1][134] <= 18'h0002c;\
    linear1_weight_array[1][135] <= 18'h2007d;\
    linear1_weight_array[1][136] <= 18'h20087;\
    linear1_weight_array[1][137] <= 18'h20054;\
    linear1_weight_array[1][138] <= 18'h2005d;\
    linear1_weight_array[1][139] <= 18'h20004;\
    linear1_weight_array[1][140] <= 18'h20059;\
    linear1_weight_array[1][141] <= 18'h00026;\
    linear1_weight_array[1][142] <= 18'h2001d;\
    linear1_weight_array[1][143] <= 18'h2004d;\
    linear1_weight_array[1][144] <= 18'h0003f;\
    linear1_weight_array[1][145] <= 18'h2003b;\
    linear1_weight_array[1][146] <= 18'h2004c;\
    linear1_weight_array[1][147] <= 18'h20074;\
    linear1_weight_array[1][148] <= 18'h0000b;\
    linear1_weight_array[1][149] <= 18'h20019;\
    linear1_weight_array[2][0] <= 18'h000c8;\
    linear1_weight_array[2][1] <= 18'h2005d;\
    linear1_weight_array[2][2] <= 18'h20095;\
    linear1_weight_array[2][3] <= 18'h20038;\
    linear1_weight_array[2][4] <= 18'h0008d;\
    linear1_weight_array[2][5] <= 18'h00159;\
    linear1_weight_array[2][6] <= 18'h0008b;\
    linear1_weight_array[2][7] <= 18'h2006d;\
    linear1_weight_array[2][8] <= 18'h000a7;\
    linear1_weight_array[2][9] <= 18'h20088;\
    linear1_weight_array[2][10] <= 18'h00249;\
    linear1_weight_array[2][11] <= 18'h00070;\
    linear1_weight_array[2][12] <= 18'h00095;\
    linear1_weight_array[2][13] <= 18'h000ef;\
    linear1_weight_array[2][14] <= 18'h001d1;\
    linear1_weight_array[2][15] <= 18'h00099;\
    linear1_weight_array[2][16] <= 18'h2007b;\
    linear1_weight_array[2][17] <= 18'h200b7;\
    linear1_weight_array[2][18] <= 18'h20051;\
    linear1_weight_array[2][19] <= 18'h00167;\
    linear1_weight_array[2][20] <= 18'h200f1;\
    linear1_weight_array[2][21] <= 18'h200ba;\
    linear1_weight_array[2][22] <= 18'h20087;\
    linear1_weight_array[2][23] <= 18'h20039;\
    linear1_weight_array[2][24] <= 18'h0002d;\
    linear1_weight_array[2][25] <= 18'h00055;\
    linear1_weight_array[2][26] <= 18'h0003f;\
    linear1_weight_array[2][27] <= 18'h0016a;\
    linear1_weight_array[2][28] <= 18'h0003e;\
    linear1_weight_array[2][29] <= 18'h20152;\
    linear1_weight_array[2][30] <= 18'h200c1;\
    linear1_weight_array[2][31] <= 18'h2012a;\
    linear1_weight_array[2][32] <= 18'h200b8;\
    linear1_weight_array[2][33] <= 18'h2007f;\
    linear1_weight_array[2][34] <= 18'h20150;\
    linear1_weight_array[2][35] <= 18'h2015e;\
    linear1_weight_array[2][36] <= 18'h20053;\
    linear1_weight_array[2][37] <= 18'h2000e;\
    linear1_weight_array[2][38] <= 18'h201b9;\
    linear1_weight_array[2][39] <= 18'h00124;\
    linear1_weight_array[2][40] <= 18'h2000d;\
    linear1_weight_array[2][41] <= 18'h00130;\
    linear1_weight_array[2][42] <= 18'h00125;\
    linear1_weight_array[2][43] <= 18'h000a9;\
    linear1_weight_array[2][44] <= 18'h20003;\
    linear1_weight_array[2][45] <= 18'h000ff;\
    linear1_weight_array[2][46] <= 18'h000da;\
    linear1_weight_array[2][47] <= 18'h0004e;\
    linear1_weight_array[2][48] <= 18'h201ac;\
    linear1_weight_array[2][49] <= 18'h200fd;\
    linear1_weight_array[2][50] <= 18'h0045d;\
    linear1_weight_array[2][51] <= 18'h000d2;\
    linear1_weight_array[2][52] <= 18'h000d8;\
    linear1_weight_array[2][53] <= 18'h000eb;\
    linear1_weight_array[2][54] <= 18'h00128;\
    linear1_weight_array[2][55] <= 18'h20135;\
    linear1_weight_array[2][56] <= 18'h200be;\
    linear1_weight_array[2][57] <= 18'h2000b;\
    linear1_weight_array[2][58] <= 18'h000aa;\
    linear1_weight_array[2][59] <= 18'h20030;\
    linear1_weight_array[2][60] <= 18'h20033;\
    linear1_weight_array[2][61] <= 18'h201c8;\
    linear1_weight_array[2][62] <= 18'h00071;\
    linear1_weight_array[2][63] <= 18'h000f6;\
    linear1_weight_array[2][64] <= 18'h2005b;\
    linear1_weight_array[2][65] <= 18'h0045d;\
    linear1_weight_array[2][66] <= 18'h00037;\
    linear1_weight_array[2][67] <= 18'h00021;\
    linear1_weight_array[2][68] <= 18'h00079;\
    linear1_weight_array[2][69] <= 18'h20061;\
    linear1_weight_array[2][70] <= 18'h00236;\
    linear1_weight_array[2][71] <= 18'h20170;\
    linear1_weight_array[2][72] <= 18'h20045;\
    linear1_weight_array[2][73] <= 18'h2002a;\
    linear1_weight_array[2][74] <= 18'h20023;\
    linear1_weight_array[2][75] <= 18'h00035;\
    linear1_weight_array[2][76] <= 18'h20112;\
    linear1_weight_array[2][77] <= 18'h2003a;\
    linear1_weight_array[2][78] <= 18'h00051;\
    linear1_weight_array[2][79] <= 18'h0009b;\
    linear1_weight_array[2][80] <= 18'h20009;\
    linear1_weight_array[2][81] <= 18'h200b4;\
    linear1_weight_array[2][82] <= 18'h20006;\
    linear1_weight_array[2][83] <= 18'h00150;\
    linear1_weight_array[2][84] <= 18'h001c1;\
    linear1_weight_array[2][85] <= 18'h00112;\
    linear1_weight_array[2][86] <= 18'h0003f;\
    linear1_weight_array[2][87] <= 18'h0007a;\
    linear1_weight_array[2][88] <= 18'h00002;\
    linear1_weight_array[2][89] <= 18'h00083;\
    linear1_weight_array[2][90] <= 18'h000ce;\
    linear1_weight_array[2][91] <= 18'h0015c;\
    linear1_weight_array[2][92] <= 18'h000b5;\
    linear1_weight_array[2][93] <= 18'h00021;\
    linear1_weight_array[2][94] <= 18'h2009f;\
    linear1_weight_array[2][95] <= 18'h200a5;\
    linear1_weight_array[2][96] <= 18'h00087;\
    linear1_weight_array[2][97] <= 18'h0001b;\
    linear1_weight_array[2][98] <= 18'h00048;\
    linear1_weight_array[2][99] <= 18'h20180;\
    linear1_weight_array[2][100] <= 18'h00128;\
    linear1_weight_array[2][101] <= 18'h000c4;\
    linear1_weight_array[2][102] <= 18'h000d6;\
    linear1_weight_array[2][103] <= 18'h20053;\
    linear1_weight_array[2][104] <= 18'h20157;\
    linear1_weight_array[2][105] <= 18'h200aa;\
    linear1_weight_array[2][106] <= 18'h200f2;\
    linear1_weight_array[2][107] <= 18'h20056;\
    linear1_weight_array[2][108] <= 18'h20068;\
    linear1_weight_array[2][109] <= 18'h201ff;\
    linear1_weight_array[2][110] <= 18'h200e0;\
    linear1_weight_array[2][111] <= 18'h20101;\
    linear1_weight_array[2][112] <= 18'h000d7;\
    linear1_weight_array[2][113] <= 18'h00114;\
    linear1_weight_array[2][114] <= 18'h0003d;\
    linear1_weight_array[2][115] <= 18'h20041;\
    linear1_weight_array[2][116] <= 18'h20065;\
    linear1_weight_array[2][117] <= 18'h0004f;\
    linear1_weight_array[2][118] <= 18'h0017d;\
    linear1_weight_array[2][119] <= 18'h20000;\
    linear1_weight_array[2][120] <= 18'h000f4;\
    linear1_weight_array[2][121] <= 18'h00029;\
    linear1_weight_array[2][122] <= 18'h20044;\
    linear1_weight_array[2][123] <= 18'h000ef;\
    linear1_weight_array[2][124] <= 18'h000f2;\
    linear1_weight_array[2][125] <= 18'h000ea;\
    linear1_weight_array[2][126] <= 18'h0011d;\
    linear1_weight_array[2][127] <= 18'h00033;\
    linear1_weight_array[2][128] <= 18'h200c4;\
    linear1_weight_array[2][129] <= 18'h20273;\
    linear1_weight_array[2][130] <= 18'h00226;\
    linear1_weight_array[2][131] <= 18'h0001c;\
    linear1_weight_array[2][132] <= 18'h00024;\
    linear1_weight_array[2][133] <= 18'h00000;\
    linear1_weight_array[2][134] <= 18'h000a7;\
    linear1_weight_array[2][135] <= 18'h0002d;\
    linear1_weight_array[2][136] <= 18'h200a2;\
    linear1_weight_array[2][137] <= 18'h00056;\
    linear1_weight_array[2][138] <= 18'h00014;\
    linear1_weight_array[2][139] <= 18'h2002d;\
    linear1_weight_array[2][140] <= 18'h200c4;\
    linear1_weight_array[2][141] <= 18'h00013;\
    linear1_weight_array[2][142] <= 18'h000dd;\
    linear1_weight_array[2][143] <= 18'h0004e;\
    linear1_weight_array[2][144] <= 18'h0016a;\
    linear1_weight_array[2][145] <= 18'h2001f;\
    linear1_weight_array[2][146] <= 18'h00083;\
    linear1_weight_array[2][147] <= 18'h00055;\
    linear1_weight_array[2][148] <= 18'h00090;\
    linear1_weight_array[2][149] <= 18'h0009f;\
    linear1_weight_array[3][0] <= 18'h2007d;\
    linear1_weight_array[3][1] <= 18'h20081;\
    linear1_weight_array[3][2] <= 18'h20051;\
    linear1_weight_array[3][3] <= 18'h00024;\
    linear1_weight_array[3][4] <= 18'h0001f;\
    linear1_weight_array[3][5] <= 18'h20110;\
    linear1_weight_array[3][6] <= 18'h2004b;\
    linear1_weight_array[3][7] <= 18'h00111;\
    linear1_weight_array[3][8] <= 18'h0011c;\
    linear1_weight_array[3][9] <= 18'h20101;\
    linear1_weight_array[3][10] <= 18'h20206;\
    linear1_weight_array[3][11] <= 18'h2015b;\
    linear1_weight_array[3][12] <= 18'h20021;\
    linear1_weight_array[3][13] <= 18'h00075;\
    linear1_weight_array[3][14] <= 18'h0002b;\
    linear1_weight_array[3][15] <= 18'h203cb;\
    linear1_weight_array[3][16] <= 18'h000a7;\
    linear1_weight_array[3][17] <= 18'h200a9;\
    linear1_weight_array[3][18] <= 18'h2001a;\
    linear1_weight_array[3][19] <= 18'h20206;\
    linear1_weight_array[3][20] <= 18'h200de;\
    linear1_weight_array[3][21] <= 18'h00034;\
    linear1_weight_array[3][22] <= 18'h000e4;\
    linear1_weight_array[3][23] <= 18'h20215;\
    linear1_weight_array[3][24] <= 18'h20209;\
    linear1_weight_array[3][25] <= 18'h2001a;\
    linear1_weight_array[3][26] <= 18'h20146;\
    linear1_weight_array[3][27] <= 18'h200d2;\
    linear1_weight_array[3][28] <= 18'h0006f;\
    linear1_weight_array[3][29] <= 18'h000b3;\
    linear1_weight_array[3][30] <= 18'h200d4;\
    linear1_weight_array[3][31] <= 18'h2015b;\
    linear1_weight_array[3][32] <= 18'h200e8;\
    linear1_weight_array[3][33] <= 18'h00090;\
    linear1_weight_array[3][34] <= 18'h001f2;\
    linear1_weight_array[3][35] <= 18'h00088;\
    linear1_weight_array[3][36] <= 18'h2008a;\
    linear1_weight_array[3][37] <= 18'h200ba;\
    linear1_weight_array[3][38] <= 18'h00029;\
    linear1_weight_array[3][39] <= 18'h00063;\
    linear1_weight_array[3][40] <= 18'h000d9;\
    linear1_weight_array[3][41] <= 18'h000ed;\
    linear1_weight_array[3][42] <= 18'h20018;\
    linear1_weight_array[3][43] <= 18'h20132;\
    linear1_weight_array[3][44] <= 18'h202e7;\
    linear1_weight_array[3][45] <= 18'h20019;\
    linear1_weight_array[3][46] <= 18'h000a2;\
    linear1_weight_array[3][47] <= 18'h000bc;\
    linear1_weight_array[3][48] <= 18'h2004b;\
    linear1_weight_array[3][49] <= 18'h20152;\
    linear1_weight_array[3][50] <= 18'h00061;\
    linear1_weight_array[3][51] <= 18'h001a8;\
    linear1_weight_array[3][52] <= 18'h00083;\
    linear1_weight_array[3][53] <= 18'h20021;\
    linear1_weight_array[3][54] <= 18'h20020;\
    linear1_weight_array[3][55] <= 18'h000ea;\
    linear1_weight_array[3][56] <= 18'h00099;\
    linear1_weight_array[3][57] <= 18'h00157;\
    linear1_weight_array[3][58] <= 18'h20082;\
    linear1_weight_array[3][59] <= 18'h200ea;\
    linear1_weight_array[3][60] <= 18'h00070;\
    linear1_weight_array[3][61] <= 18'h00071;\
    linear1_weight_array[3][62] <= 18'h20045;\
    linear1_weight_array[3][63] <= 18'h200be;\
    linear1_weight_array[3][64] <= 18'h000d8;\
    linear1_weight_array[3][65] <= 18'h0022d;\
    linear1_weight_array[3][66] <= 18'h000ac;\
    linear1_weight_array[3][67] <= 18'h200dd;\
    linear1_weight_array[3][68] <= 18'h00003;\
    linear1_weight_array[3][69] <= 18'h00072;\
    linear1_weight_array[3][70] <= 18'h00280;\
    linear1_weight_array[3][71] <= 18'h2000d;\
    linear1_weight_array[3][72] <= 18'h20004;\
    linear1_weight_array[3][73] <= 18'h000a9;\
    linear1_weight_array[3][74] <= 18'h2007f;\
    linear1_weight_array[3][75] <= 18'h2001c;\
    linear1_weight_array[3][76] <= 18'h200a0;\
    linear1_weight_array[3][77] <= 18'h000e1;\
    linear1_weight_array[3][78] <= 18'h00139;\
    linear1_weight_array[3][79] <= 18'h0001b;\
    linear1_weight_array[3][80] <= 18'h20030;\
    linear1_weight_array[3][81] <= 18'h000b8;\
    linear1_weight_array[3][82] <= 18'h00063;\
    linear1_weight_array[3][83] <= 18'h2002a;\
    linear1_weight_array[3][84] <= 18'h2004c;\
    linear1_weight_array[3][85] <= 18'h000c6;\
    linear1_weight_array[3][86] <= 18'h00118;\
    linear1_weight_array[3][87] <= 18'h200e2;\
    linear1_weight_array[3][88] <= 18'h2009b;\
    linear1_weight_array[3][89] <= 18'h000eb;\
    linear1_weight_array[3][90] <= 18'h2009e;\
    linear1_weight_array[3][91] <= 18'h000da;\
    linear1_weight_array[3][92] <= 18'h00002;\
    linear1_weight_array[3][93] <= 18'h000d8;\
    linear1_weight_array[3][94] <= 18'h0008e;\
    linear1_weight_array[3][95] <= 18'h20070;\
    linear1_weight_array[3][96] <= 18'h00036;\
    linear1_weight_array[3][97] <= 18'h200c4;\
    linear1_weight_array[3][98] <= 18'h00144;\
    linear1_weight_array[3][99] <= 18'h001a0;\
    linear1_weight_array[3][100] <= 18'h00060;\
    linear1_weight_array[3][101] <= 18'h202af;\
    linear1_weight_array[3][102] <= 18'h20026;\
    linear1_weight_array[3][103] <= 18'h00136;\
    linear1_weight_array[3][104] <= 18'h0008d;\
    linear1_weight_array[3][105] <= 18'h20194;\
    linear1_weight_array[3][106] <= 18'h20154;\
    linear1_weight_array[3][107] <= 18'h2002b;\
    linear1_weight_array[3][108] <= 18'h0001a;\
    linear1_weight_array[3][109] <= 18'h00199;\
    linear1_weight_array[3][110] <= 18'h2000f;\
    linear1_weight_array[3][111] <= 18'h00049;\
    linear1_weight_array[3][112] <= 18'h200a4;\
    linear1_weight_array[3][113] <= 18'h20083;\
    linear1_weight_array[3][114] <= 18'h0003b;\
    linear1_weight_array[3][115] <= 18'h000d3;\
    linear1_weight_array[3][116] <= 18'h000ec;\
    linear1_weight_array[3][117] <= 18'h00076;\
    linear1_weight_array[3][118] <= 18'h000df;\
    linear1_weight_array[3][119] <= 18'h200ab;\
    linear1_weight_array[3][120] <= 18'h0002e;\
    linear1_weight_array[3][121] <= 18'h20043;\
    linear1_weight_array[3][122] <= 18'h00046;\
    linear1_weight_array[3][123] <= 18'h00080;\
    linear1_weight_array[3][124] <= 18'h0004f;\
    linear1_weight_array[3][125] <= 18'h0001b;\
    linear1_weight_array[3][126] <= 18'h00025;\
    linear1_weight_array[3][127] <= 18'h2010e;\
    linear1_weight_array[3][128] <= 18'h00036;\
    linear1_weight_array[3][129] <= 18'h00037;\
    linear1_weight_array[3][130] <= 18'h2015c;\
    linear1_weight_array[3][131] <= 18'h2009a;\
    linear1_weight_array[3][132] <= 18'h2004e;\
    linear1_weight_array[3][133] <= 18'h20084;\
    linear1_weight_array[3][134] <= 18'h202ba;\
    linear1_weight_array[3][135] <= 18'h20262;\
    linear1_weight_array[3][136] <= 18'h20057;\
    linear1_weight_array[3][137] <= 18'h2007f;\
    linear1_weight_array[3][138] <= 18'h20027;\
    linear1_weight_array[3][139] <= 18'h000e6;\
    linear1_weight_array[3][140] <= 18'h0009e;\
    linear1_weight_array[3][141] <= 18'h00020;\
    linear1_weight_array[3][142] <= 18'h00007;\
    linear1_weight_array[3][143] <= 18'h00190;\
    linear1_weight_array[3][144] <= 18'h00104;\
    linear1_weight_array[3][145] <= 18'h0007c;\
    linear1_weight_array[3][146] <= 18'h000c4;\
    linear1_weight_array[3][147] <= 18'h0006d;\
    linear1_weight_array[3][148] <= 18'h00046;\
    linear1_weight_array[3][149] <= 18'h000bf;\
    linear1_weight_array[4][0] <= 18'h2003f;\
    linear1_weight_array[4][1] <= 18'h2002d;\
    linear1_weight_array[4][2] <= 18'h00028;\
    linear1_weight_array[4][3] <= 18'h00033;\
    linear1_weight_array[4][4] <= 18'h0001d;\
    linear1_weight_array[4][5] <= 18'h2005f;\
    linear1_weight_array[4][6] <= 18'h00018;\
    linear1_weight_array[4][7] <= 18'h2001c;\
    linear1_weight_array[4][8] <= 18'h20028;\
    linear1_weight_array[4][9] <= 18'h0000c;\
    linear1_weight_array[4][10] <= 18'h20064;\
    linear1_weight_array[4][11] <= 18'h20037;\
    linear1_weight_array[4][12] <= 18'h2000b;\
    linear1_weight_array[4][13] <= 18'h2001d;\
    linear1_weight_array[4][14] <= 18'h20051;\
    linear1_weight_array[4][15] <= 18'h00010;\
    linear1_weight_array[4][16] <= 18'h2004c;\
    linear1_weight_array[4][17] <= 18'h20046;\
    linear1_weight_array[4][18] <= 18'h0004c;\
    linear1_weight_array[4][19] <= 18'h20049;\
    linear1_weight_array[4][20] <= 18'h20059;\
    linear1_weight_array[4][21] <= 18'h00008;\
    linear1_weight_array[4][22] <= 18'h00018;\
    linear1_weight_array[4][23] <= 18'h20001;\
    linear1_weight_array[4][24] <= 18'h00023;\
    linear1_weight_array[4][25] <= 18'h20003;\
    linear1_weight_array[4][26] <= 18'h2000e;\
    linear1_weight_array[4][27] <= 18'h20007;\
    linear1_weight_array[4][28] <= 18'h20009;\
    linear1_weight_array[4][29] <= 18'h2001d;\
    linear1_weight_array[4][30] <= 18'h2000f;\
    linear1_weight_array[4][31] <= 18'h20034;\
    linear1_weight_array[4][32] <= 18'h20018;\
    linear1_weight_array[4][33] <= 18'h0004f;\
    linear1_weight_array[4][34] <= 18'h0001c;\
    linear1_weight_array[4][35] <= 18'h2001d;\
    linear1_weight_array[4][36] <= 18'h20069;\
    linear1_weight_array[4][37] <= 18'h20066;\
    linear1_weight_array[4][38] <= 18'h20022;\
    linear1_weight_array[4][39] <= 18'h20052;\
    linear1_weight_array[4][40] <= 18'h20027;\
    linear1_weight_array[4][41] <= 18'h0002e;\
    linear1_weight_array[4][42] <= 18'h0001d;\
    linear1_weight_array[4][43] <= 18'h00007;\
    linear1_weight_array[4][44] <= 18'h00018;\
    linear1_weight_array[4][45] <= 18'h20062;\
    linear1_weight_array[4][46] <= 18'h2003a;\
    linear1_weight_array[4][47] <= 18'h00023;\
    linear1_weight_array[4][48] <= 18'h0000d;\
    linear1_weight_array[4][49] <= 18'h00032;\
    linear1_weight_array[4][50] <= 18'h0001d;\
    linear1_weight_array[4][51] <= 18'h0001e;\
    linear1_weight_array[4][52] <= 18'h20003;\
    linear1_weight_array[4][53] <= 18'h00000;\
    linear1_weight_array[4][54] <= 18'h0000d;\
    linear1_weight_array[4][55] <= 18'h00025;\
    linear1_weight_array[4][56] <= 18'h20012;\
    linear1_weight_array[4][57] <= 18'h20022;\
    linear1_weight_array[4][58] <= 18'h00035;\
    linear1_weight_array[4][59] <= 18'h0000f;\
    linear1_weight_array[4][60] <= 18'h2001c;\
    linear1_weight_array[4][61] <= 18'h20043;\
    linear1_weight_array[4][62] <= 18'h0003f;\
    linear1_weight_array[4][63] <= 18'h00000;\
    linear1_weight_array[4][64] <= 18'h20056;\
    linear1_weight_array[4][65] <= 18'h0000a;\
    linear1_weight_array[4][66] <= 18'h2002a;\
    linear1_weight_array[4][67] <= 18'h0002d;\
    linear1_weight_array[4][68] <= 18'h00007;\
    linear1_weight_array[4][69] <= 18'h2005d;\
    linear1_weight_array[4][70] <= 18'h20031;\
    linear1_weight_array[4][71] <= 18'h2005c;\
    linear1_weight_array[4][72] <= 18'h20054;\
    linear1_weight_array[4][73] <= 18'h20053;\
    linear1_weight_array[4][74] <= 18'h2003c;\
    linear1_weight_array[4][75] <= 18'h20028;\
    linear1_weight_array[4][76] <= 18'h20049;\
    linear1_weight_array[4][77] <= 18'h20039;\
    linear1_weight_array[4][78] <= 18'h2000a;\
    linear1_weight_array[4][79] <= 18'h20066;\
    linear1_weight_array[4][80] <= 18'h2003c;\
    linear1_weight_array[4][81] <= 18'h20040;\
    linear1_weight_array[4][82] <= 18'h20017;\
    linear1_weight_array[4][83] <= 18'h20033;\
    linear1_weight_array[4][84] <= 18'h2003f;\
    linear1_weight_array[4][85] <= 18'h2000d;\
    linear1_weight_array[4][86] <= 18'h20042;\
    linear1_weight_array[4][87] <= 18'h20062;\
    linear1_weight_array[4][88] <= 18'h20065;\
    linear1_weight_array[4][89] <= 18'h2006a;\
    linear1_weight_array[4][90] <= 18'h20006;\
    linear1_weight_array[4][91] <= 18'h20020;\
    linear1_weight_array[4][92] <= 18'h2004b;\
    linear1_weight_array[4][93] <= 18'h20045;\
    linear1_weight_array[4][94] <= 18'h20026;\
    linear1_weight_array[4][95] <= 18'h2003c;\
    linear1_weight_array[4][96] <= 18'h20061;\
    linear1_weight_array[4][97] <= 18'h00008;\
    linear1_weight_array[4][98] <= 18'h2004a;\
    linear1_weight_array[4][99] <= 18'h20003;\
    linear1_weight_array[4][100] <= 18'h00010;\
    linear1_weight_array[4][101] <= 18'h00054;\
    linear1_weight_array[4][102] <= 18'h20018;\
    linear1_weight_array[4][103] <= 18'h00027;\
    linear1_weight_array[4][104] <= 18'h20054;\
    linear1_weight_array[4][105] <= 18'h2006d;\
    linear1_weight_array[4][106] <= 18'h0003a;\
    linear1_weight_array[4][107] <= 18'h00001;\
    linear1_weight_array[4][108] <= 18'h20043;\
    linear1_weight_array[4][109] <= 18'h2003f;\
    linear1_weight_array[4][110] <= 18'h20013;\
    linear1_weight_array[4][111] <= 18'h2002a;\
    linear1_weight_array[4][112] <= 18'h20009;\
    linear1_weight_array[4][113] <= 18'h20061;\
    linear1_weight_array[4][114] <= 18'h0005e;\
    linear1_weight_array[4][115] <= 18'h0001f;\
    linear1_weight_array[4][116] <= 18'h0000e;\
    linear1_weight_array[4][117] <= 18'h20059;\
    linear1_weight_array[4][118] <= 18'h00000;\
    linear1_weight_array[4][119] <= 18'h00007;\
    linear1_weight_array[4][120] <= 18'h00030;\
    linear1_weight_array[4][121] <= 18'h00035;\
    linear1_weight_array[4][122] <= 18'h2005d;\
    linear1_weight_array[4][123] <= 18'h00014;\
    linear1_weight_array[4][124] <= 18'h00000;\
    linear1_weight_array[4][125] <= 18'h0002b;\
    linear1_weight_array[4][126] <= 18'h2000a;\
    linear1_weight_array[4][127] <= 18'h2001b;\
    linear1_weight_array[4][128] <= 18'h20015;\
    linear1_weight_array[4][129] <= 18'h20041;\
    linear1_weight_array[4][130] <= 18'h0000d;\
    linear1_weight_array[4][131] <= 18'h0003a;\
    linear1_weight_array[4][132] <= 18'h2003b;\
    linear1_weight_array[4][133] <= 18'h00005;\
    linear1_weight_array[4][134] <= 18'h00018;\
    linear1_weight_array[4][135] <= 18'h20003;\
    linear1_weight_array[4][136] <= 18'h20011;\
    linear1_weight_array[4][137] <= 18'h20021;\
    linear1_weight_array[4][138] <= 18'h0000a;\
    linear1_weight_array[4][139] <= 18'h2003d;\
    linear1_weight_array[4][140] <= 18'h2006c;\
    linear1_weight_array[4][141] <= 18'h20039;\
    linear1_weight_array[4][142] <= 18'h0000b;\
    linear1_weight_array[4][143] <= 18'h20078;\
    linear1_weight_array[4][144] <= 18'h20012;\
    linear1_weight_array[4][145] <= 18'h2004a;\
    linear1_weight_array[4][146] <= 18'h20027;\
    linear1_weight_array[4][147] <= 18'h00003;\
    linear1_weight_array[4][148] <= 18'h20055;\
    linear1_weight_array[4][149] <= 18'h2001b;\
    linear1_weight_array[5][0] <= 18'h20000;\
    linear1_weight_array[5][1] <= 18'h20063;\
    linear1_weight_array[5][2] <= 18'h2007a;\
    linear1_weight_array[5][3] <= 18'h20080;\
    linear1_weight_array[5][4] <= 18'h20030;\
    linear1_weight_array[5][5] <= 18'h20063;\
    linear1_weight_array[5][6] <= 18'h2009c;\
    linear1_weight_array[5][7] <= 18'h2007d;\
    linear1_weight_array[5][8] <= 18'h20029;\
    linear1_weight_array[5][9] <= 18'h00048;\
    linear1_weight_array[5][10] <= 18'h0000e;\
    linear1_weight_array[5][11] <= 18'h2005e;\
    linear1_weight_array[5][12] <= 18'h00066;\
    linear1_weight_array[5][13] <= 18'h00083;\
    linear1_weight_array[5][14] <= 18'h00173;\
    linear1_weight_array[5][15] <= 18'h00207;\
    linear1_weight_array[5][16] <= 18'h2003a;\
    linear1_weight_array[5][17] <= 18'h00011;\
    linear1_weight_array[5][18] <= 18'h00081;\
    linear1_weight_array[5][19] <= 18'h000ed;\
    linear1_weight_array[5][20] <= 18'h00128;\
    linear1_weight_array[5][21] <= 18'h00067;\
    linear1_weight_array[5][22] <= 18'h2004b;\
    linear1_weight_array[5][23] <= 18'h00035;\
    linear1_weight_array[5][24] <= 18'h20165;\
    linear1_weight_array[5][25] <= 18'h0000a;\
    linear1_weight_array[5][26] <= 18'h000dc;\
    linear1_weight_array[5][27] <= 18'h200a0;\
    linear1_weight_array[5][28] <= 18'h201b6;\
    linear1_weight_array[5][29] <= 18'h200cd;\
    linear1_weight_array[5][30] <= 18'h00043;\
    linear1_weight_array[5][31] <= 18'h20043;\
    linear1_weight_array[5][32] <= 18'h20115;\
    linear1_weight_array[5][33] <= 18'h2013f;\
    linear1_weight_array[5][34] <= 18'h0014e;\
    linear1_weight_array[5][35] <= 18'h0011c;\
    linear1_weight_array[5][36] <= 18'h00230;\
    linear1_weight_array[5][37] <= 18'h000ac;\
    linear1_weight_array[5][38] <= 18'h20016;\
    linear1_weight_array[5][39] <= 18'h00013;\
    linear1_weight_array[5][40] <= 18'h2007b;\
    linear1_weight_array[5][41] <= 18'h000c6;\
    linear1_weight_array[5][42] <= 18'h0008f;\
    linear1_weight_array[5][43] <= 18'h000c9;\
    linear1_weight_array[5][44] <= 18'h000a9;\
    linear1_weight_array[5][45] <= 18'h00109;\
    linear1_weight_array[5][46] <= 18'h200ef;\
    linear1_weight_array[5][47] <= 18'h20098;\
    linear1_weight_array[5][48] <= 18'h20030;\
    linear1_weight_array[5][49] <= 18'h0016f;\
    linear1_weight_array[5][50] <= 18'h2009d;\
    linear1_weight_array[5][51] <= 18'h0010e;\
    linear1_weight_array[5][52] <= 18'h000b8;\
    linear1_weight_array[5][53] <= 18'h00114;\
    linear1_weight_array[5][54] <= 18'h00142;\
    linear1_weight_array[5][55] <= 18'h00173;\
    linear1_weight_array[5][56] <= 18'h000b1;\
    linear1_weight_array[5][57] <= 18'h20013;\
    linear1_weight_array[5][58] <= 18'h2004d;\
    linear1_weight_array[5][59] <= 18'h20039;\
    linear1_weight_array[5][60] <= 18'h20082;\
    linear1_weight_array[5][61] <= 18'h00019;\
    linear1_weight_array[5][62] <= 18'h00007;\
    linear1_weight_array[5][63] <= 18'h200b4;\
    linear1_weight_array[5][64] <= 18'h200b5;\
    linear1_weight_array[5][65] <= 18'h201a1;\
    linear1_weight_array[5][66] <= 18'h20255;\
    linear1_weight_array[5][67] <= 18'h200d9;\
    linear1_weight_array[5][68] <= 18'h00027;\
    linear1_weight_array[5][69] <= 18'h0005e;\
    linear1_weight_array[5][70] <= 18'h20131;\
    linear1_weight_array[5][71] <= 18'h200d7;\
    linear1_weight_array[5][72] <= 18'h000e6;\
    linear1_weight_array[5][73] <= 18'h0007f;\
    linear1_weight_array[5][74] <= 18'h00154;\
    linear1_weight_array[5][75] <= 18'h200a2;\
    linear1_weight_array[5][76] <= 18'h200cc;\
    linear1_weight_array[5][77] <= 18'h200a5;\
    linear1_weight_array[5][78] <= 18'h20057;\
    linear1_weight_array[5][79] <= 18'h00137;\
    linear1_weight_array[5][80] <= 18'h2008d;\
    linear1_weight_array[5][81] <= 18'h00079;\
    linear1_weight_array[5][82] <= 18'h0014e;\
    linear1_weight_array[5][83] <= 18'h00046;\
    linear1_weight_array[5][84] <= 18'h20039;\
    linear1_weight_array[5][85] <= 18'h000c3;\
    linear1_weight_array[5][86] <= 18'h0007f;\
    linear1_weight_array[5][87] <= 18'h00050;\
    linear1_weight_array[5][88] <= 18'h2010e;\
    linear1_weight_array[5][89] <= 18'h20127;\
    linear1_weight_array[5][90] <= 18'h200ad;\
    linear1_weight_array[5][91] <= 18'h200a9;\
    linear1_weight_array[5][92] <= 18'h2001e;\
    linear1_weight_array[5][93] <= 18'h00043;\
    linear1_weight_array[5][94] <= 18'h000ba;\
    linear1_weight_array[5][95] <= 18'h000bd;\
    linear1_weight_array[5][96] <= 18'h20084;\
    linear1_weight_array[5][97] <= 18'h000dc;\
    linear1_weight_array[5][98] <= 18'h20015;\
    linear1_weight_array[5][99] <= 18'h001bc;\
    linear1_weight_array[5][100] <= 18'h0017c;\
    linear1_weight_array[5][101] <= 18'h00031;\
    linear1_weight_array[5][102] <= 18'h200ed;\
    linear1_weight_array[5][103] <= 18'h0000f;\
    linear1_weight_array[5][104] <= 18'h20054;\
    linear1_weight_array[5][105] <= 18'h00124;\
    linear1_weight_array[5][106] <= 18'h00004;\
    linear1_weight_array[5][107] <= 18'h20037;\
    linear1_weight_array[5][108] <= 18'h2001d;\
    linear1_weight_array[5][109] <= 18'h2005a;\
    linear1_weight_array[5][110] <= 18'h000b1;\
    linear1_weight_array[5][111] <= 18'h0011c;\
    linear1_weight_array[5][112] <= 18'h000dc;\
    linear1_weight_array[5][113] <= 18'h0009e;\
    linear1_weight_array[5][114] <= 18'h200ea;\
    linear1_weight_array[5][115] <= 18'h2000e;\
    linear1_weight_array[5][116] <= 18'h00037;\
    linear1_weight_array[5][117] <= 18'h00062;\
    linear1_weight_array[5][118] <= 18'h200a3;\
    linear1_weight_array[5][119] <= 18'h200bb;\
    linear1_weight_array[5][120] <= 18'h200a5;\
    linear1_weight_array[5][121] <= 18'h2006a;\
    linear1_weight_array[5][122] <= 18'h2001d;\
    linear1_weight_array[5][123] <= 18'h200e1;\
    linear1_weight_array[5][124] <= 18'h20072;\
    linear1_weight_array[5][125] <= 18'h00047;\
    linear1_weight_array[5][126] <= 18'h0002c;\
    linear1_weight_array[5][127] <= 18'h00080;\
    linear1_weight_array[5][128] <= 18'h000dc;\
    linear1_weight_array[5][129] <= 18'h002d5;\
    linear1_weight_array[5][130] <= 18'h20042;\
    linear1_weight_array[5][131] <= 18'h0001c;\
    linear1_weight_array[5][132] <= 18'h000e1;\
    linear1_weight_array[5][133] <= 18'h200d0;\
    linear1_weight_array[5][134] <= 18'h003c9;\
    linear1_weight_array[5][135] <= 18'h0012d;\
    linear1_weight_array[5][136] <= 18'h000c3;\
    linear1_weight_array[5][137] <= 18'h00139;\
    linear1_weight_array[5][138] <= 18'h00077;\
    linear1_weight_array[5][139] <= 18'h20215;\
    linear1_weight_array[5][140] <= 18'h00121;\
    linear1_weight_array[5][141] <= 18'h00020;\
    linear1_weight_array[5][142] <= 18'h0006c;\
    linear1_weight_array[5][143] <= 18'h20059;\
    linear1_weight_array[5][144] <= 18'h20182;\
    linear1_weight_array[5][145] <= 18'h0006b;\
    linear1_weight_array[5][146] <= 18'h00013;\
    linear1_weight_array[5][147] <= 18'h0006a;\
    linear1_weight_array[5][148] <= 18'h00082;\
    linear1_weight_array[5][149] <= 18'h20044;\
    linear1_weight_array[6][0] <= 18'h00068;\
    linear1_weight_array[6][1] <= 18'h000af;\
    linear1_weight_array[6][2] <= 18'h0006d;\
    linear1_weight_array[6][3] <= 18'h00068;\
    linear1_weight_array[6][4] <= 18'h0000a;\
    linear1_weight_array[6][5] <= 18'h0015f;\
    linear1_weight_array[6][6] <= 18'h000be;\
    linear1_weight_array[6][7] <= 18'h0009d;\
    linear1_weight_array[6][8] <= 18'h00095;\
    linear1_weight_array[6][9] <= 18'h200d9;\
    linear1_weight_array[6][10] <= 18'h20070;\
    linear1_weight_array[6][11] <= 18'h20078;\
    linear1_weight_array[6][12] <= 18'h2005f;\
    linear1_weight_array[6][13] <= 18'h000b6;\
    linear1_weight_array[6][14] <= 18'h0003b;\
    linear1_weight_array[6][15] <= 18'h2001a;\
    linear1_weight_array[6][16] <= 18'h2001e;\
    linear1_weight_array[6][17] <= 18'h00081;\
    linear1_weight_array[6][18] <= 18'h2000f;\
    linear1_weight_array[6][19] <= 18'h000c7;\
    linear1_weight_array[6][20] <= 18'h001dd;\
    linear1_weight_array[6][21] <= 18'h20044;\
    linear1_weight_array[6][22] <= 18'h000c6;\
    linear1_weight_array[6][23] <= 18'h00104;\
    linear1_weight_array[6][24] <= 18'h200dd;\
    linear1_weight_array[6][25] <= 18'h20004;\
    linear1_weight_array[6][26] <= 18'h00083;\
    linear1_weight_array[6][27] <= 18'h0008c;\
    linear1_weight_array[6][28] <= 18'h00003;\
    linear1_weight_array[6][29] <= 18'h2012c;\
    linear1_weight_array[6][30] <= 18'h0003b;\
    linear1_weight_array[6][31] <= 18'h200fd;\
    linear1_weight_array[6][32] <= 18'h20002;\
    linear1_weight_array[6][33] <= 18'h20003;\
    linear1_weight_array[6][34] <= 18'h20118;\
    linear1_weight_array[6][35] <= 18'h20063;\
    linear1_weight_array[6][36] <= 18'h20042;\
    linear1_weight_array[6][37] <= 18'h00001;\
    linear1_weight_array[6][38] <= 18'h201ee;\
    linear1_weight_array[6][39] <= 18'h2014e;\
    linear1_weight_array[6][40] <= 18'h00080;\
    linear1_weight_array[6][41] <= 18'h0002f;\
    linear1_weight_array[6][42] <= 18'h00028;\
    linear1_weight_array[6][43] <= 18'h00044;\
    linear1_weight_array[6][44] <= 18'h201ee;\
    linear1_weight_array[6][45] <= 18'h20144;\
    linear1_weight_array[6][46] <= 18'h2004b;\
    linear1_weight_array[6][47] <= 18'h00052;\
    linear1_weight_array[6][48] <= 18'h001cc;\
    linear1_weight_array[6][49] <= 18'h2004b;\
    linear1_weight_array[6][50] <= 18'h20056;\
    linear1_weight_array[6][51] <= 18'h20112;\
    linear1_weight_array[6][52] <= 18'h000b2;\
    linear1_weight_array[6][53] <= 18'h0006b;\
    linear1_weight_array[6][54] <= 18'h00107;\
    linear1_weight_array[6][55] <= 18'h20106;\
    linear1_weight_array[6][56] <= 18'h00184;\
    linear1_weight_array[6][57] <= 18'h20112;\
    linear1_weight_array[6][58] <= 18'h000f3;\
    linear1_weight_array[6][59] <= 18'h000af;\
    linear1_weight_array[6][60] <= 18'h000d7;\
    linear1_weight_array[6][61] <= 18'h000eb;\
    linear1_weight_array[6][62] <= 18'h20038;\
    linear1_weight_array[6][63] <= 18'h00021;\
    linear1_weight_array[6][64] <= 18'h00061;\
    linear1_weight_array[6][65] <= 18'h20021;\
    linear1_weight_array[6][66] <= 18'h20027;\
    linear1_weight_array[6][67] <= 18'h20019;\
    linear1_weight_array[6][68] <= 18'h000e4;\
    linear1_weight_array[6][69] <= 18'h000b9;\
    linear1_weight_array[6][70] <= 18'h20117;\
    linear1_weight_array[6][71] <= 18'h00167;\
    linear1_weight_array[6][72] <= 18'h000fe;\
    linear1_weight_array[6][73] <= 18'h0011d;\
    linear1_weight_array[6][74] <= 18'h0010b;\
    linear1_weight_array[6][75] <= 18'h2003d;\
    linear1_weight_array[6][76] <= 18'h20008;\
    linear1_weight_array[6][77] <= 18'h00003;\
    linear1_weight_array[6][78] <= 18'h00050;\
    linear1_weight_array[6][79] <= 18'h20046;\
    linear1_weight_array[6][80] <= 18'h20061;\
    linear1_weight_array[6][81] <= 18'h20008;\
    linear1_weight_array[6][82] <= 18'h000aa;\
    linear1_weight_array[6][83] <= 18'h00070;\
    linear1_weight_array[6][84] <= 18'h20012;\
    linear1_weight_array[6][85] <= 18'h20191;\
    linear1_weight_array[6][86] <= 18'h20084;\
    linear1_weight_array[6][87] <= 18'h000a4;\
    linear1_weight_array[6][88] <= 18'h0004a;\
    linear1_weight_array[6][89] <= 18'h00118;\
    linear1_weight_array[6][90] <= 18'h20081;\
    linear1_weight_array[6][91] <= 18'h20195;\
    linear1_weight_array[6][92] <= 18'h000c9;\
    linear1_weight_array[6][93] <= 18'h000ca;\
    linear1_weight_array[6][94] <= 18'h001f8;\
    linear1_weight_array[6][95] <= 18'h0016f;\
    linear1_weight_array[6][96] <= 18'h20076;\
    linear1_weight_array[6][97] <= 18'h00093;\
    linear1_weight_array[6][98] <= 18'h20021;\
    linear1_weight_array[6][99] <= 18'h201d4;\
    linear1_weight_array[6][100] <= 18'h00209;\
    linear1_weight_array[6][101] <= 18'h0014b;\
    linear1_weight_array[6][102] <= 18'h00027;\
    linear1_weight_array[6][103] <= 18'h00056;\
    linear1_weight_array[6][104] <= 18'h2003c;\
    linear1_weight_array[6][105] <= 18'h0004b;\
    linear1_weight_array[6][106] <= 18'h00043;\
    linear1_weight_array[6][107] <= 18'h20098;\
    linear1_weight_array[6][108] <= 18'h00007;\
    linear1_weight_array[6][109] <= 18'h00060;\
    linear1_weight_array[6][110] <= 18'h2006d;\
    linear1_weight_array[6][111] <= 18'h00001;\
    linear1_weight_array[6][112] <= 18'h20042;\
    linear1_weight_array[6][113] <= 18'h000b0;\
    linear1_weight_array[6][114] <= 18'h20015;\
    linear1_weight_array[6][115] <= 18'h20099;\
    linear1_weight_array[6][116] <= 18'h0003d;\
    linear1_weight_array[6][117] <= 18'h20145;\
    linear1_weight_array[6][118] <= 18'h201f5;\
    linear1_weight_array[6][119] <= 18'h200fa;\
    linear1_weight_array[6][120] <= 18'h20122;\
    linear1_weight_array[6][121] <= 18'h20060;\
    linear1_weight_array[6][122] <= 18'h2018d;\
    linear1_weight_array[6][123] <= 18'h2008d;\
    linear1_weight_array[6][124] <= 18'h20046;\
    linear1_weight_array[6][125] <= 18'h00119;\
    linear1_weight_array[6][126] <= 18'h00161;\
    linear1_weight_array[6][127] <= 18'h000db;\
    linear1_weight_array[6][128] <= 18'h2009e;\
    linear1_weight_array[6][129] <= 18'h00030;\
    linear1_weight_array[6][130] <= 18'h0003b;\
    linear1_weight_array[6][131] <= 18'h000ac;\
    linear1_weight_array[6][132] <= 18'h00027;\
    linear1_weight_array[6][133] <= 18'h0000c;\
    linear1_weight_array[6][134] <= 18'h0010e;\
    linear1_weight_array[6][135] <= 18'h00153;\
    linear1_weight_array[6][136] <= 18'h0011c;\
    linear1_weight_array[6][137] <= 18'h00185;\
    linear1_weight_array[6][138] <= 18'h0002f;\
    linear1_weight_array[6][139] <= 18'h0001a;\
    linear1_weight_array[6][140] <= 18'h00111;\
    linear1_weight_array[6][141] <= 18'h2006e;\
    linear1_weight_array[6][142] <= 18'h20048;\
    linear1_weight_array[6][143] <= 18'h20026;\
    linear1_weight_array[6][144] <= 18'h00095;\
    linear1_weight_array[6][145] <= 18'h20083;\
    linear1_weight_array[6][146] <= 18'h20116;\
    linear1_weight_array[6][147] <= 18'h20103;\
    linear1_weight_array[6][148] <= 18'h20138;\
    linear1_weight_array[6][149] <= 18'h200fe;\
    linear1_weight_array[7][0] <= 18'h00011;\
    linear1_weight_array[7][1] <= 18'h2000e;\
    linear1_weight_array[7][2] <= 18'h00046;\
    linear1_weight_array[7][3] <= 18'h000b5;\
    linear1_weight_array[7][4] <= 18'h20018;\
    linear1_weight_array[7][5] <= 18'h2009a;\
    linear1_weight_array[7][6] <= 18'h20068;\
    linear1_weight_array[7][7] <= 18'h2011a;\
    linear1_weight_array[7][8] <= 18'h20088;\
    linear1_weight_array[7][9] <= 18'h00028;\
    linear1_weight_array[7][10] <= 18'h20075;\
    linear1_weight_array[7][11] <= 18'h000ae;\
    linear1_weight_array[7][12] <= 18'h00063;\
    linear1_weight_array[7][13] <= 18'h20000;\
    linear1_weight_array[7][14] <= 18'h0002a;\
    linear1_weight_array[7][15] <= 18'h20234;\
    linear1_weight_array[7][16] <= 18'h200e1;\
    linear1_weight_array[7][17] <= 18'h0012a;\
    linear1_weight_array[7][18] <= 18'h000d7;\
    linear1_weight_array[7][19] <= 18'h0005d;\
    linear1_weight_array[7][20] <= 18'h201fb;\
    linear1_weight_array[7][21] <= 18'h200d9;\
    linear1_weight_array[7][22] <= 18'h00030;\
    linear1_weight_array[7][23] <= 18'h20029;\
    linear1_weight_array[7][24] <= 18'h00240;\
    linear1_weight_array[7][25] <= 18'h2007e;\
    linear1_weight_array[7][26] <= 18'h2000e;\
    linear1_weight_array[7][27] <= 18'h20001;\
    linear1_weight_array[7][28] <= 18'h00201;\
    linear1_weight_array[7][29] <= 18'h00009;\
    linear1_weight_array[7][30] <= 18'h000b3;\
    linear1_weight_array[7][31] <= 18'h00114;\
    linear1_weight_array[7][32] <= 18'h20017;\
    linear1_weight_array[7][33] <= 18'h00001;\
    linear1_weight_array[7][34] <= 18'h200db;\
    linear1_weight_array[7][35] <= 18'h20001;\
    linear1_weight_array[7][36] <= 18'h0004b;\
    linear1_weight_array[7][37] <= 18'h20092;\
    linear1_weight_array[7][38] <= 18'h0005b;\
    linear1_weight_array[7][39] <= 18'h0000f;\
    linear1_weight_array[7][40] <= 18'h00011;\
    linear1_weight_array[7][41] <= 18'h20065;\
    linear1_weight_array[7][42] <= 18'h2007a;\
    linear1_weight_array[7][43] <= 18'h000d1;\
    linear1_weight_array[7][44] <= 18'h2003b;\
    linear1_weight_array[7][45] <= 18'h20115;\
    linear1_weight_array[7][46] <= 18'h0001a;\
    linear1_weight_array[7][47] <= 18'h00006;\
    linear1_weight_array[7][48] <= 18'h00109;\
    linear1_weight_array[7][49] <= 18'h0000c;\
    linear1_weight_array[7][50] <= 18'h201f7;\
    linear1_weight_array[7][51] <= 18'h00005;\
    linear1_weight_array[7][52] <= 18'h0004e;\
    linear1_weight_array[7][53] <= 18'h00022;\
    linear1_weight_array[7][54] <= 18'h000e0;\
    linear1_weight_array[7][55] <= 18'h20027;\
    linear1_weight_array[7][56] <= 18'h00057;\
    linear1_weight_array[7][57] <= 18'h201da;\
    linear1_weight_array[7][58] <= 18'h00054;\
    linear1_weight_array[7][59] <= 18'h0016d;\
    linear1_weight_array[7][60] <= 18'h0000c;\
    linear1_weight_array[7][61] <= 18'h00008;\
    linear1_weight_array[7][62] <= 18'h00070;\
    linear1_weight_array[7][63] <= 18'h0006f;\
    linear1_weight_array[7][64] <= 18'h0002a;\
    linear1_weight_array[7][65] <= 18'h2011a;\
    linear1_weight_array[7][66] <= 18'h00033;\
    linear1_weight_array[7][67] <= 18'h00090;\
    linear1_weight_array[7][68] <= 18'h20006;\
    linear1_weight_array[7][69] <= 18'h20088;\
    linear1_weight_array[7][70] <= 18'h20044;\
    linear1_weight_array[7][71] <= 18'h20065;\
    linear1_weight_array[7][72] <= 18'h20076;\
    linear1_weight_array[7][73] <= 18'h20074;\
    linear1_weight_array[7][74] <= 18'h000cd;\
    linear1_weight_array[7][75] <= 18'h0004d;\
    linear1_weight_array[7][76] <= 18'h0006d;\
    linear1_weight_array[7][77] <= 18'h200fa;\
    linear1_weight_array[7][78] <= 18'h20141;\
    linear1_weight_array[7][79] <= 18'h00099;\
    linear1_weight_array[7][80] <= 18'h000d2;\
    linear1_weight_array[7][81] <= 18'h00020;\
    linear1_weight_array[7][82] <= 18'h20042;\
    linear1_weight_array[7][83] <= 18'h20042;\
    linear1_weight_array[7][84] <= 18'h0025b;\
    linear1_weight_array[7][85] <= 18'h000c1;\
    linear1_weight_array[7][86] <= 18'h000b7;\
    linear1_weight_array[7][87] <= 18'h0015e;\
    linear1_weight_array[7][88] <= 18'h0028a;\
    linear1_weight_array[7][89] <= 18'h20013;\
    linear1_weight_array[7][90] <= 18'h0010a;\
    linear1_weight_array[7][91] <= 18'h00177;\
    linear1_weight_array[7][92] <= 18'h000b1;\
    linear1_weight_array[7][93] <= 18'h20067;\
    linear1_weight_array[7][94] <= 18'h00017;\
    linear1_weight_array[7][95] <= 18'h200f1;\
    linear1_weight_array[7][96] <= 18'h20031;\
    linear1_weight_array[7][97] <= 18'h20085;\
    linear1_weight_array[7][98] <= 18'h200df;\
    linear1_weight_array[7][99] <= 18'h201c4;\
    linear1_weight_array[7][100] <= 18'h201a4;\
    linear1_weight_array[7][101] <= 18'h2000a;\
    linear1_weight_array[7][102] <= 18'h20027;\
    linear1_weight_array[7][103] <= 18'h00174;\
    linear1_weight_array[7][104] <= 18'h000dc;\
    linear1_weight_array[7][105] <= 18'h000f2;\
    linear1_weight_array[7][106] <= 18'h0018a;\
    linear1_weight_array[7][107] <= 18'h000d6;\
    linear1_weight_array[7][108] <= 18'h2010d;\
    linear1_weight_array[7][109] <= 18'h20011;\
    linear1_weight_array[7][110] <= 18'h000aa;\
    linear1_weight_array[7][111] <= 18'h00171;\
    linear1_weight_array[7][112] <= 18'h00088;\
    linear1_weight_array[7][113] <= 18'h200cd;\
    linear1_weight_array[7][114] <= 18'h20002;\
    linear1_weight_array[7][115] <= 18'h000b2;\
    linear1_weight_array[7][116] <= 18'h00052;\
    linear1_weight_array[7][117] <= 18'h20079;\
    linear1_weight_array[7][118] <= 18'h200d9;\
    linear1_weight_array[7][119] <= 18'h000c1;\
    linear1_weight_array[7][120] <= 18'h001a3;\
    linear1_weight_array[7][121] <= 18'h00139;\
    linear1_weight_array[7][122] <= 18'h000a9;\
    linear1_weight_array[7][123] <= 18'h00094;\
    linear1_weight_array[7][124] <= 18'h00153;\
    linear1_weight_array[7][125] <= 18'h00027;\
    linear1_weight_array[7][126] <= 18'h200cd;\
    linear1_weight_array[7][127] <= 18'h200ba;\
    linear1_weight_array[7][128] <= 18'h200af;\
    linear1_weight_array[7][129] <= 18'h20097;\
    linear1_weight_array[7][130] <= 18'h201e4;\
    linear1_weight_array[7][131] <= 18'h200b8;\
    linear1_weight_array[7][132] <= 18'h00007;\
    linear1_weight_array[7][133] <= 18'h000b2;\
    linear1_weight_array[7][134] <= 18'h200de;\
    linear1_weight_array[7][135] <= 18'h2002b;\
    linear1_weight_array[7][136] <= 18'h2001d;\
    linear1_weight_array[7][137] <= 18'h0009b;\
    linear1_weight_array[7][138] <= 18'h0012f;\
    linear1_weight_array[7][139] <= 18'h00112;\
    linear1_weight_array[7][140] <= 18'h2006e;\
    linear1_weight_array[7][141] <= 18'h00036;\
    linear1_weight_array[7][142] <= 18'h2003b;\
    linear1_weight_array[7][143] <= 18'h2007a;\
    linear1_weight_array[7][144] <= 18'h0002a;\
    linear1_weight_array[7][145] <= 18'h20043;\
    linear1_weight_array[7][146] <= 18'h20078;\
    linear1_weight_array[7][147] <= 18'h20078;\
    linear1_weight_array[7][148] <= 18'h20028;\
    linear1_weight_array[7][149] <= 18'h20047;\
    linear1_weight_array[8][0] <= 18'h20010;\
    linear1_weight_array[8][1] <= 18'h0001f;\
    linear1_weight_array[8][2] <= 18'h00028;\
    linear1_weight_array[8][3] <= 18'h00016;\
    linear1_weight_array[8][4] <= 18'h2001f;\
    linear1_weight_array[8][5] <= 18'h00009;\
    linear1_weight_array[8][6] <= 18'h00015;\
    linear1_weight_array[8][7] <= 18'h20002;\
    linear1_weight_array[8][8] <= 18'h2004f;\
    linear1_weight_array[8][9] <= 18'h2001d;\
    linear1_weight_array[8][10] <= 18'h00033;\
    linear1_weight_array[8][11] <= 18'h20036;\
    linear1_weight_array[8][12] <= 18'h20058;\
    linear1_weight_array[8][13] <= 18'h0000a;\
    linear1_weight_array[8][14] <= 18'h00022;\
    linear1_weight_array[8][15] <= 18'h20000;\
    linear1_weight_array[8][16] <= 18'h2002d;\
    linear1_weight_array[8][17] <= 18'h00008;\
    linear1_weight_array[8][18] <= 18'h00000;\
    linear1_weight_array[8][19] <= 18'h20018;\
    linear1_weight_array[8][20] <= 18'h0002c;\
    linear1_weight_array[8][21] <= 18'h00023;\
    linear1_weight_array[8][22] <= 18'h0003d;\
    linear1_weight_array[8][23] <= 18'h00014;\
    linear1_weight_array[8][24] <= 18'h00021;\
    linear1_weight_array[8][25] <= 18'h20023;\
    linear1_weight_array[8][26] <= 18'h20032;\
    linear1_weight_array[8][27] <= 18'h20057;\
    linear1_weight_array[8][28] <= 18'h20054;\
    linear1_weight_array[8][29] <= 18'h00014;\
    linear1_weight_array[8][30] <= 18'h00021;\
    linear1_weight_array[8][31] <= 18'h00038;\
    linear1_weight_array[8][32] <= 18'h20044;\
    linear1_weight_array[8][33] <= 18'h20044;\
    linear1_weight_array[8][34] <= 18'h2001d;\
    linear1_weight_array[8][35] <= 18'h20036;\
    linear1_weight_array[8][36] <= 18'h20059;\
    linear1_weight_array[8][37] <= 18'h20054;\
    linear1_weight_array[8][38] <= 18'h0001d;\
    linear1_weight_array[8][39] <= 18'h20036;\
    linear1_weight_array[8][40] <= 18'h00000;\
    linear1_weight_array[8][41] <= 18'h00005;\
    linear1_weight_array[8][42] <= 18'h20054;\
    linear1_weight_array[8][43] <= 18'h20036;\
    linear1_weight_array[8][44] <= 18'h20021;\
    linear1_weight_array[8][45] <= 18'h2001d;\
    linear1_weight_array[8][46] <= 18'h2001e;\
    linear1_weight_array[8][47] <= 18'h00010;\
    linear1_weight_array[8][48] <= 18'h2005d;\
    linear1_weight_array[8][49] <= 18'h00004;\
    linear1_weight_array[8][50] <= 18'h20005;\
    linear1_weight_array[8][51] <= 18'h00015;\
    linear1_weight_array[8][52] <= 18'h20038;\
    linear1_weight_array[8][53] <= 18'h00010;\
    linear1_weight_array[8][54] <= 18'h20036;\
    linear1_weight_array[8][55] <= 18'h00037;\
    linear1_weight_array[8][56] <= 18'h20044;\
    linear1_weight_array[8][57] <= 18'h00044;\
    linear1_weight_array[8][58] <= 18'h00038;\
    linear1_weight_array[8][59] <= 18'h20047;\
    linear1_weight_array[8][60] <= 18'h20043;\
    linear1_weight_array[8][61] <= 18'h20027;\
    linear1_weight_array[8][62] <= 18'h2001f;\
    linear1_weight_array[8][63] <= 18'h20040;\
    linear1_weight_array[8][64] <= 18'h0002e;\
    linear1_weight_array[8][65] <= 18'h20005;\
    linear1_weight_array[8][66] <= 18'h00051;\
    linear1_weight_array[8][67] <= 18'h20004;\
    linear1_weight_array[8][68] <= 18'h20009;\
    linear1_weight_array[8][69] <= 18'h2001d;\
    linear1_weight_array[8][70] <= 18'h2005c;\
    linear1_weight_array[8][71] <= 18'h20038;\
    linear1_weight_array[8][72] <= 18'h2001a;\
    linear1_weight_array[8][73] <= 18'h2003b;\
    linear1_weight_array[8][74] <= 18'h00015;\
    linear1_weight_array[8][75] <= 18'h0003e;\
    linear1_weight_array[8][76] <= 18'h20021;\
    linear1_weight_array[8][77] <= 18'h00012;\
    linear1_weight_array[8][78] <= 18'h2000b;\
    linear1_weight_array[8][79] <= 18'h20021;\
    linear1_weight_array[8][80] <= 18'h20029;\
    linear1_weight_array[8][81] <= 18'h20022;\
    linear1_weight_array[8][82] <= 18'h00023;\
    linear1_weight_array[8][83] <= 18'h20064;\
    linear1_weight_array[8][84] <= 18'h00016;\
    linear1_weight_array[8][85] <= 18'h00015;\
    linear1_weight_array[8][86] <= 18'h2005a;\
    linear1_weight_array[8][87] <= 18'h20023;\
    linear1_weight_array[8][88] <= 18'h0003b;\
    linear1_weight_array[8][89] <= 18'h2002f;\
    linear1_weight_array[8][90] <= 18'h20048;\
    linear1_weight_array[8][91] <= 18'h20012;\
    linear1_weight_array[8][92] <= 18'h20001;\
    linear1_weight_array[8][93] <= 18'h20052;\
    linear1_weight_array[8][94] <= 18'h20049;\
    linear1_weight_array[8][95] <= 18'h0003b;\
    linear1_weight_array[8][96] <= 18'h20015;\
    linear1_weight_array[8][97] <= 18'h20002;\
    linear1_weight_array[8][98] <= 18'h20014;\
    linear1_weight_array[8][99] <= 18'h2005c;\
    linear1_weight_array[8][100] <= 18'h00009;\
    linear1_weight_array[8][101] <= 18'h20016;\
    linear1_weight_array[8][102] <= 18'h20054;\
    linear1_weight_array[8][103] <= 18'h00037;\
    linear1_weight_array[8][104] <= 18'h00002;\
    linear1_weight_array[8][105] <= 18'h2000f;\
    linear1_weight_array[8][106] <= 18'h20011;\
    linear1_weight_array[8][107] <= 18'h20063;\
    linear1_weight_array[8][108] <= 18'h20053;\
    linear1_weight_array[8][109] <= 18'h20026;\
    linear1_weight_array[8][110] <= 18'h00026;\
    linear1_weight_array[8][111] <= 18'h0001d;\
    linear1_weight_array[8][112] <= 18'h0000c;\
    linear1_weight_array[8][113] <= 18'h0001b;\
    linear1_weight_array[8][114] <= 18'h20007;\
    linear1_weight_array[8][115] <= 18'h20066;\
    linear1_weight_array[8][116] <= 18'h20042;\
    linear1_weight_array[8][117] <= 18'h00037;\
    linear1_weight_array[8][118] <= 18'h00021;\
    linear1_weight_array[8][119] <= 18'h0001e;\
    linear1_weight_array[8][120] <= 18'h00020;\
    linear1_weight_array[8][121] <= 18'h00027;\
    linear1_weight_array[8][122] <= 18'h20003;\
    linear1_weight_array[8][123] <= 18'h2002b;\
    linear1_weight_array[8][124] <= 18'h2003b;\
    linear1_weight_array[8][125] <= 18'h20006;\
    linear1_weight_array[8][126] <= 18'h2002e;\
    linear1_weight_array[8][127] <= 18'h20008;\
    linear1_weight_array[8][128] <= 18'h2004d;\
    linear1_weight_array[8][129] <= 18'h00014;\
    linear1_weight_array[8][130] <= 18'h20005;\
    linear1_weight_array[8][131] <= 18'h20017;\
    linear1_weight_array[8][132] <= 18'h20050;\
    linear1_weight_array[8][133] <= 18'h20003;\
    linear1_weight_array[8][134] <= 18'h2000e;\
    linear1_weight_array[8][135] <= 18'h2003c;\
    linear1_weight_array[8][136] <= 18'h20023;\
    linear1_weight_array[8][137] <= 18'h2005c;\
    linear1_weight_array[8][138] <= 18'h2005c;\
    linear1_weight_array[8][139] <= 18'h20050;\
    linear1_weight_array[8][140] <= 18'h00025;\
    linear1_weight_array[8][141] <= 18'h00004;\
    linear1_weight_array[8][142] <= 18'h2004e;\
    linear1_weight_array[8][143] <= 18'h0003d;\
    linear1_weight_array[8][144] <= 18'h20062;\
    linear1_weight_array[8][145] <= 18'h0000a;\
    linear1_weight_array[8][146] <= 18'h2001e;\
    linear1_weight_array[8][147] <= 18'h0001e;\
    linear1_weight_array[8][148] <= 18'h2001b;\
    linear1_weight_array[8][149] <= 18'h0000d;\
    linear1_weight_array[9][0] <= 18'h0009d;\
    linear1_weight_array[9][1] <= 18'h00159;\
    linear1_weight_array[9][2] <= 18'h0005f;\
    linear1_weight_array[9][3] <= 18'h0002e;\
    linear1_weight_array[9][4] <= 18'h000b8;\
    linear1_weight_array[9][5] <= 18'h20115;\
    linear1_weight_array[9][6] <= 18'h000c0;\
    linear1_weight_array[9][7] <= 18'h00042;\
    linear1_weight_array[9][8] <= 18'h00008;\
    linear1_weight_array[9][9] <= 18'h0001b;\
    linear1_weight_array[9][10] <= 18'h20124;\
    linear1_weight_array[9][11] <= 18'h20163;\
    linear1_weight_array[9][12] <= 18'h2016d;\
    linear1_weight_array[9][13] <= 18'h2012d;\
    linear1_weight_array[9][14] <= 18'h201a1;\
    linear1_weight_array[9][15] <= 18'h2021b;\
    linear1_weight_array[9][16] <= 18'h00002;\
    linear1_weight_array[9][17] <= 18'h2008a;\
    linear1_weight_array[9][18] <= 18'h200fd;\
    linear1_weight_array[9][19] <= 18'h200f2;\
    linear1_weight_array[9][20] <= 18'h20019;\
    linear1_weight_array[9][21] <= 18'h00007;\
    linear1_weight_array[9][22] <= 18'h20189;\
    linear1_weight_array[9][23] <= 18'h20118;\
    linear1_weight_array[9][24] <= 18'h2014d;\
    linear1_weight_array[9][25] <= 18'h200b9;\
    linear1_weight_array[9][26] <= 18'h000c3;\
    linear1_weight_array[9][27] <= 18'h00013;\
    linear1_weight_array[9][28] <= 18'h00071;\
    linear1_weight_array[9][29] <= 18'h2004a;\
    linear1_weight_array[9][30] <= 18'h2009a;\
    linear1_weight_array[9][31] <= 18'h000a9;\
    linear1_weight_array[9][32] <= 18'h20006;\
    linear1_weight_array[9][33] <= 18'h20050;\
    linear1_weight_array[9][34] <= 18'h200ce;\
    linear1_weight_array[9][35] <= 18'h00019;\
    linear1_weight_array[9][36] <= 18'h000a8;\
    linear1_weight_array[9][37] <= 18'h000c2;\
    linear1_weight_array[9][38] <= 18'h000ee;\
    linear1_weight_array[9][39] <= 18'h20158;\
    linear1_weight_array[9][40] <= 18'h2000f;\
    linear1_weight_array[9][41] <= 18'h20067;\
    linear1_weight_array[9][42] <= 18'h00000;\
    linear1_weight_array[9][43] <= 18'h2000a;\
    linear1_weight_array[9][44] <= 18'h001c3;\
    linear1_weight_array[9][45] <= 18'h00086;\
    linear1_weight_array[9][46] <= 18'h00029;\
    linear1_weight_array[9][47] <= 18'h00011;\
    linear1_weight_array[9][48] <= 18'h20115;\
    linear1_weight_array[9][49] <= 18'h200bf;\
    linear1_weight_array[9][50] <= 18'h201cd;\
    linear1_weight_array[9][51] <= 18'h2010f;\
    linear1_weight_array[9][52] <= 18'h20070;\
    linear1_weight_array[9][53] <= 18'h0006f;\
    linear1_weight_array[9][54] <= 18'h20029;\
    linear1_weight_array[9][55] <= 18'h201d5;\
    linear1_weight_array[9][56] <= 18'h20092;\
    linear1_weight_array[9][57] <= 18'h200cb;\
    linear1_weight_array[9][58] <= 18'h00130;\
    linear1_weight_array[9][59] <= 18'h0002c;\
    linear1_weight_array[9][60] <= 18'h00032;\
    linear1_weight_array[9][61] <= 18'h00071;\
    linear1_weight_array[9][62] <= 18'h00093;\
    linear1_weight_array[9][63] <= 18'h000a0;\
    linear1_weight_array[9][64] <= 18'h20045;\
    linear1_weight_array[9][65] <= 18'h2019d;\
    linear1_weight_array[9][66] <= 18'h000ee;\
    linear1_weight_array[9][67] <= 18'h20070;\
    linear1_weight_array[9][68] <= 18'h2004c;\
    linear1_weight_array[9][69] <= 18'h2000d;\
    linear1_weight_array[9][70] <= 18'h200d8;\
    linear1_weight_array[9][71] <= 18'h20152;\
    linear1_weight_array[9][72] <= 18'h00026;\
    linear1_weight_array[9][73] <= 18'h2001b;\
    linear1_weight_array[9][74] <= 18'h20045;\
    linear1_weight_array[9][75] <= 18'h20015;\
    linear1_weight_array[9][76] <= 18'h00085;\
    linear1_weight_array[9][77] <= 18'h000a8;\
    linear1_weight_array[9][78] <= 18'h0008e;\
    linear1_weight_array[9][79] <= 18'h2013c;\
    linear1_weight_array[9][80] <= 18'h00046;\
    linear1_weight_array[9][81] <= 18'h2000e;\
    linear1_weight_array[9][82] <= 18'h00104;\
    linear1_weight_array[9][83] <= 18'h00100;\
    linear1_weight_array[9][84] <= 18'h2005d;\
    linear1_weight_array[9][85] <= 18'h200d4;\
    linear1_weight_array[9][86] <= 18'h000a2;\
    linear1_weight_array[9][87] <= 18'h00165;\
    linear1_weight_array[9][88] <= 18'h20174;\
    linear1_weight_array[9][89] <= 18'h0007c;\
    linear1_weight_array[9][90] <= 18'h00090;\
    linear1_weight_array[9][91] <= 18'h20041;\
    linear1_weight_array[9][92] <= 18'h20060;\
    linear1_weight_array[9][93] <= 18'h20119;\
    linear1_weight_array[9][94] <= 18'h20093;\
    linear1_weight_array[9][95] <= 18'h20002;\
    linear1_weight_array[9][96] <= 18'h20047;\
    linear1_weight_array[9][97] <= 18'h00066;\
    linear1_weight_array[9][98] <= 18'h00042;\
    linear1_weight_array[9][99] <= 18'h0021f;\
    linear1_weight_array[9][100] <= 18'h20045;\
    linear1_weight_array[9][101] <= 18'h200c4;\
    linear1_weight_array[9][102] <= 18'h20078;\
    linear1_weight_array[9][103] <= 18'h0006e;\
    linear1_weight_array[9][104] <= 18'h200cc;\
    linear1_weight_array[9][105] <= 18'h000ec;\
    linear1_weight_array[9][106] <= 18'h0010b;\
    linear1_weight_array[9][107] <= 18'h0002a;\
    linear1_weight_array[9][108] <= 18'h200ef;\
    linear1_weight_array[9][109] <= 18'h20178;\
    linear1_weight_array[9][110] <= 18'h000db;\
    linear1_weight_array[9][111] <= 18'h0013c;\
    linear1_weight_array[9][112] <= 18'h000af;\
    linear1_weight_array[9][113] <= 18'h001fb;\
    linear1_weight_array[9][114] <= 18'h00026;\
    linear1_weight_array[9][115] <= 18'h2003b;\
    linear1_weight_array[9][116] <= 18'h00076;\
    linear1_weight_array[9][117] <= 18'h000e0;\
    linear1_weight_array[9][118] <= 18'h00008;\
    linear1_weight_array[9][119] <= 18'h20379;\
    linear1_weight_array[9][120] <= 18'h00178;\
    linear1_weight_array[9][121] <= 18'h0001e;\
    linear1_weight_array[9][122] <= 18'h2007e;\
    linear1_weight_array[9][123] <= 18'h00093;\
    linear1_weight_array[9][124] <= 18'h2005b;\
    linear1_weight_array[9][125] <= 18'h0007f;\
    linear1_weight_array[9][126] <= 18'h00002;\
    linear1_weight_array[9][127] <= 18'h2006d;\
    linear1_weight_array[9][128] <= 18'h2007f;\
    linear1_weight_array[9][129] <= 18'h20128;\
    linear1_weight_array[9][130] <= 18'h2006a;\
    linear1_weight_array[9][131] <= 18'h200c3;\
    linear1_weight_array[9][132] <= 18'h20025;\
    linear1_weight_array[9][133] <= 18'h20096;\
    linear1_weight_array[9][134] <= 18'h2007e;\
    linear1_weight_array[9][135] <= 18'h200fa;\
    linear1_weight_array[9][136] <= 18'h00029;\
    linear1_weight_array[9][137] <= 18'h00093;\
    linear1_weight_array[9][138] <= 18'h000b3;\
    linear1_weight_array[9][139] <= 18'h00026;\
    linear1_weight_array[9][140] <= 18'h200d6;\
    linear1_weight_array[9][141] <= 18'h2000f;\
    linear1_weight_array[9][142] <= 18'h00049;\
    linear1_weight_array[9][143] <= 18'h20110;\
    linear1_weight_array[9][144] <= 18'h200a0;\
    linear1_weight_array[9][145] <= 18'h00002;\
    linear1_weight_array[9][146] <= 18'h000b7;\
    linear1_weight_array[9][147] <= 18'h00076;\
    linear1_weight_array[9][148] <= 18'h0011f;\
    linear1_weight_array[9][149] <= 18'h00019;\
    linear1_weight_array[10][0] <= 18'h20039;\
    linear1_weight_array[10][1] <= 18'h00004;\
    linear1_weight_array[10][2] <= 18'h2005b;\
    linear1_weight_array[10][3] <= 18'h20058;\
    linear1_weight_array[10][4] <= 18'h20022;\
    linear1_weight_array[10][5] <= 18'h20012;\
    linear1_weight_array[10][6] <= 18'h0001d;\
    linear1_weight_array[10][7] <= 18'h20031;\
    linear1_weight_array[10][8] <= 18'h0001b;\
    linear1_weight_array[10][9] <= 18'h0002d;\
    linear1_weight_array[10][10] <= 18'h20005;\
    linear1_weight_array[10][11] <= 18'h2002f;\
    linear1_weight_array[10][12] <= 18'h20016;\
    linear1_weight_array[10][13] <= 18'h20019;\
    linear1_weight_array[10][14] <= 18'h2006e;\
    linear1_weight_array[10][15] <= 18'h20003;\
    linear1_weight_array[10][16] <= 18'h00028;\
    linear1_weight_array[10][17] <= 18'h20038;\
    linear1_weight_array[10][18] <= 18'h2001c;\
    linear1_weight_array[10][19] <= 18'h20051;\
    linear1_weight_array[10][20] <= 18'h20019;\
    linear1_weight_array[10][21] <= 18'h0003f;\
    linear1_weight_array[10][22] <= 18'h00013;\
    linear1_weight_array[10][23] <= 18'h20057;\
    linear1_weight_array[10][24] <= 18'h0000b;\
    linear1_weight_array[10][25] <= 18'h20075;\
    linear1_weight_array[10][26] <= 18'h00028;\
    linear1_weight_array[10][27] <= 18'h00021;\
    linear1_weight_array[10][28] <= 18'h20043;\
    linear1_weight_array[10][29] <= 18'h20081;\
    linear1_weight_array[10][30] <= 18'h2007b;\
    linear1_weight_array[10][31] <= 18'h00023;\
    linear1_weight_array[10][32] <= 18'h20001;\
    linear1_weight_array[10][33] <= 18'h00013;\
    linear1_weight_array[10][34] <= 18'h0001a;\
    linear1_weight_array[10][35] <= 18'h20017;\
    linear1_weight_array[10][36] <= 18'h2000d;\
    linear1_weight_array[10][37] <= 18'h00005;\
    linear1_weight_array[10][38] <= 18'h20018;\
    linear1_weight_array[10][39] <= 18'h0003a;\
    linear1_weight_array[10][40] <= 18'h20015;\
    linear1_weight_array[10][41] <= 18'h2003f;\
    linear1_weight_array[10][42] <= 18'h20062;\
    linear1_weight_array[10][43] <= 18'h00042;\
    linear1_weight_array[10][44] <= 18'h20052;\
    linear1_weight_array[10][45] <= 18'h20043;\
    linear1_weight_array[10][46] <= 18'h00011;\
    linear1_weight_array[10][47] <= 18'h20060;\
    linear1_weight_array[10][48] <= 18'h20003;\
    linear1_weight_array[10][49] <= 18'h2000b;\
    linear1_weight_array[10][50] <= 18'h0002a;\
    linear1_weight_array[10][51] <= 18'h0002d;\
    linear1_weight_array[10][52] <= 18'h20056;\
    linear1_weight_array[10][53] <= 18'h2007a;\
    linear1_weight_array[10][54] <= 18'h20035;\
    linear1_weight_array[10][55] <= 18'h0002c;\
    linear1_weight_array[10][56] <= 18'h2003d;\
    linear1_weight_array[10][57] <= 18'h2003d;\
    linear1_weight_array[10][58] <= 18'h20008;\
    linear1_weight_array[10][59] <= 18'h20020;\
    linear1_weight_array[10][60] <= 18'h00021;\
    linear1_weight_array[10][61] <= 18'h00026;\
    linear1_weight_array[10][62] <= 18'h00019;\
    linear1_weight_array[10][63] <= 18'h2001d;\
    linear1_weight_array[10][64] <= 18'h20025;\
    linear1_weight_array[10][65] <= 18'h2001c;\
    linear1_weight_array[10][66] <= 18'h20015;\
    linear1_weight_array[10][67] <= 18'h2003e;\
    linear1_weight_array[10][68] <= 18'h2003d;\
    linear1_weight_array[10][69] <= 18'h20056;\
    linear1_weight_array[10][70] <= 18'h2005f;\
    linear1_weight_array[10][71] <= 18'h2003e;\
    linear1_weight_array[10][72] <= 18'h00034;\
    linear1_weight_array[10][73] <= 18'h20005;\
    linear1_weight_array[10][74] <= 18'h00027;\
    linear1_weight_array[10][75] <= 18'h20069;\
    linear1_weight_array[10][76] <= 18'h20021;\
    linear1_weight_array[10][77] <= 18'h20066;\
    linear1_weight_array[10][78] <= 18'h20039;\
    linear1_weight_array[10][79] <= 18'h20054;\
    linear1_weight_array[10][80] <= 18'h00018;\
    linear1_weight_array[10][81] <= 18'h00013;\
    linear1_weight_array[10][82] <= 18'h2000c;\
    linear1_weight_array[10][83] <= 18'h20009;\
    linear1_weight_array[10][84] <= 18'h20030;\
    linear1_weight_array[10][85] <= 18'h00014;\
    linear1_weight_array[10][86] <= 18'h2005c;\
    linear1_weight_array[10][87] <= 18'h20062;\
    linear1_weight_array[10][88] <= 18'h2002a;\
    linear1_weight_array[10][89] <= 18'h2005a;\
    linear1_weight_array[10][90] <= 18'h0002b;\
    linear1_weight_array[10][91] <= 18'h0001d;\
    linear1_weight_array[10][92] <= 18'h20015;\
    linear1_weight_array[10][93] <= 18'h00007;\
    linear1_weight_array[10][94] <= 18'h0000a;\
    linear1_weight_array[10][95] <= 18'h00024;\
    linear1_weight_array[10][96] <= 18'h20041;\
    linear1_weight_array[10][97] <= 18'h2005a;\
    linear1_weight_array[10][98] <= 18'h20009;\
    linear1_weight_array[10][99] <= 18'h0000f;\
    linear1_weight_array[10][100] <= 18'h20001;\
    linear1_weight_array[10][101] <= 18'h20040;\
    linear1_weight_array[10][102] <= 18'h20033;\
    linear1_weight_array[10][103] <= 18'h20035;\
    linear1_weight_array[10][104] <= 18'h2000a;\
    linear1_weight_array[10][105] <= 18'h00018;\
    linear1_weight_array[10][106] <= 18'h20021;\
    linear1_weight_array[10][107] <= 18'h20001;\
    linear1_weight_array[10][108] <= 18'h00023;\
    linear1_weight_array[10][109] <= 18'h00020;\
    linear1_weight_array[10][110] <= 18'h2002a;\
    linear1_weight_array[10][111] <= 18'h20010;\
    linear1_weight_array[10][112] <= 18'h20006;\
    linear1_weight_array[10][113] <= 18'h2007e;\
    linear1_weight_array[10][114] <= 18'h0001c;\
    linear1_weight_array[10][115] <= 18'h20032;\
    linear1_weight_array[10][116] <= 18'h2000c;\
    linear1_weight_array[10][117] <= 18'h2003a;\
    linear1_weight_array[10][118] <= 18'h0000e;\
    linear1_weight_array[10][119] <= 18'h20012;\
    linear1_weight_array[10][120] <= 18'h20022;\
    linear1_weight_array[10][121] <= 18'h00046;\
    linear1_weight_array[10][122] <= 18'h20052;\
    linear1_weight_array[10][123] <= 18'h0001c;\
    linear1_weight_array[10][124] <= 18'h20021;\
    linear1_weight_array[10][125] <= 18'h20001;\
    linear1_weight_array[10][126] <= 18'h0001b;\
    linear1_weight_array[10][127] <= 18'h20041;\
    linear1_weight_array[10][128] <= 18'h20046;\
    linear1_weight_array[10][129] <= 18'h2000d;\
    linear1_weight_array[10][130] <= 18'h00049;\
    linear1_weight_array[10][131] <= 18'h00002;\
    linear1_weight_array[10][132] <= 18'h2002c;\
    linear1_weight_array[10][133] <= 18'h20030;\
    linear1_weight_array[10][134] <= 18'h00025;\
    linear1_weight_array[10][135] <= 18'h20022;\
    linear1_weight_array[10][136] <= 18'h20006;\
    linear1_weight_array[10][137] <= 18'h2006c;\
    linear1_weight_array[10][138] <= 18'h2001a;\
    linear1_weight_array[10][139] <= 18'h2002b;\
    linear1_weight_array[10][140] <= 18'h2000a;\
    linear1_weight_array[10][141] <= 18'h00011;\
    linear1_weight_array[10][142] <= 18'h20036;\
    linear1_weight_array[10][143] <= 18'h00030;\
    linear1_weight_array[10][144] <= 18'h2007d;\
    linear1_weight_array[10][145] <= 18'h00010;\
    linear1_weight_array[10][146] <= 18'h20007;\
    linear1_weight_array[10][147] <= 18'h00025;\
    linear1_weight_array[10][148] <= 18'h2003f;\
    linear1_weight_array[10][149] <= 18'h0003a;\
    linear1_weight_array[11][0] <= 18'h000ec;\
    linear1_weight_array[11][1] <= 18'h000f6;\
    linear1_weight_array[11][2] <= 18'h00094;\
    linear1_weight_array[11][3] <= 18'h20027;\
    linear1_weight_array[11][4] <= 18'h20056;\
    linear1_weight_array[11][5] <= 18'h00194;\
    linear1_weight_array[11][6] <= 18'h20025;\
    linear1_weight_array[11][7] <= 18'h20020;\
    linear1_weight_array[11][8] <= 18'h200ca;\
    linear1_weight_array[11][9] <= 18'h2014f;\
    linear1_weight_array[11][10] <= 18'h000a9;\
    linear1_weight_array[11][11] <= 18'h2000d;\
    linear1_weight_array[11][12] <= 18'h2009a;\
    linear1_weight_array[11][13] <= 18'h2006b;\
    linear1_weight_array[11][14] <= 18'h00073;\
    linear1_weight_array[11][15] <= 18'h0006a;\
    linear1_weight_array[11][16] <= 18'h000d8;\
    linear1_weight_array[11][17] <= 18'h00051;\
    linear1_weight_array[11][18] <= 18'h2006a;\
    linear1_weight_array[11][19] <= 18'h00068;\
    linear1_weight_array[11][20] <= 18'h0024b;\
    linear1_weight_array[11][21] <= 18'h0005e;\
    linear1_weight_array[11][22] <= 18'h00051;\
    linear1_weight_array[11][23] <= 18'h00016;\
    linear1_weight_array[11][24] <= 18'h0018c;\
    linear1_weight_array[11][25] <= 18'h00005;\
    linear1_weight_array[11][26] <= 18'h00040;\
    linear1_weight_array[11][27] <= 18'h001bc;\
    linear1_weight_array[11][28] <= 18'h00225;\
    linear1_weight_array[11][29] <= 18'h00256;\
    linear1_weight_array[11][30] <= 18'h2013a;\
    linear1_weight_array[11][31] <= 18'h20109;\
    linear1_weight_array[11][32] <= 18'h2006d;\
    linear1_weight_array[11][33] <= 18'h00021;\
    linear1_weight_array[11][34] <= 18'h200a4;\
    linear1_weight_array[11][35] <= 18'h20022;\
    linear1_weight_array[11][36] <= 18'h000f9;\
    linear1_weight_array[11][37] <= 18'h00015;\
    linear1_weight_array[11][38] <= 18'h20048;\
    linear1_weight_array[11][39] <= 18'h200a2;\
    linear1_weight_array[11][40] <= 18'h000a6;\
    linear1_weight_array[11][41] <= 18'h20045;\
    linear1_weight_array[11][42] <= 18'h20048;\
    linear1_weight_array[11][43] <= 18'h00014;\
    linear1_weight_array[11][44] <= 18'h00003;\
    linear1_weight_array[11][45] <= 18'h2005d;\
    linear1_weight_array[11][46] <= 18'h20059;\
    linear1_weight_array[11][47] <= 18'h2006e;\
    linear1_weight_array[11][48] <= 18'h0010d;\
    linear1_weight_array[11][49] <= 18'h001a7;\
    linear1_weight_array[11][50] <= 18'h20246;\
    linear1_weight_array[11][51] <= 18'h2020f;\
    linear1_weight_array[11][52] <= 18'h00040;\
    linear1_weight_array[11][53] <= 18'h2001c;\
    linear1_weight_array[11][54] <= 18'h000cf;\
    linear1_weight_array[11][55] <= 18'h0004a;\
    linear1_weight_array[11][56] <= 18'h200c6;\
    linear1_weight_array[11][57] <= 18'h200aa;\
    linear1_weight_array[11][58] <= 18'h0004d;\
    linear1_weight_array[11][59] <= 18'h00131;\
    linear1_weight_array[11][60] <= 18'h002fe;\
    linear1_weight_array[11][61] <= 18'h2010f;\
    linear1_weight_array[11][62] <= 18'h2004b;\
    linear1_weight_array[11][63] <= 18'h2005c;\
    linear1_weight_array[11][64] <= 18'h00086;\
    linear1_weight_array[11][65] <= 18'h0011c;\
    linear1_weight_array[11][66] <= 18'h20167;\
    linear1_weight_array[11][67] <= 18'h200fb;\
    linear1_weight_array[11][68] <= 18'h00015;\
    linear1_weight_array[11][69] <= 18'h00028;\
    linear1_weight_array[11][70] <= 18'h00032;\
    linear1_weight_array[11][71] <= 18'h000d8;\
    linear1_weight_array[11][72] <= 18'h00000;\
    linear1_weight_array[11][73] <= 18'h2009a;\
    linear1_weight_array[11][74] <= 18'h2001c;\
    linear1_weight_array[11][75] <= 18'h00020;\
    linear1_weight_array[11][76] <= 18'h200ae;\
    linear1_weight_array[11][77] <= 18'h2005c;\
    linear1_weight_array[11][78] <= 18'h2008d;\
    linear1_weight_array[11][79] <= 18'h0004e;\
    linear1_weight_array[11][80] <= 18'h20014;\
    linear1_weight_array[11][81] <= 18'h00002;\
    linear1_weight_array[11][82] <= 18'h00057;\
    linear1_weight_array[11][83] <= 18'h0004a;\
    linear1_weight_array[11][84] <= 18'h00006;\
    linear1_weight_array[11][85] <= 18'h00052;\
    linear1_weight_array[11][86] <= 18'h00008;\
    linear1_weight_array[11][87] <= 18'h201b7;\
    linear1_weight_array[11][88] <= 18'h000b7;\
    linear1_weight_array[11][89] <= 18'h00278;\
    linear1_weight_array[11][90] <= 18'h20063;\
    linear1_weight_array[11][91] <= 18'h20029;\
    linear1_weight_array[11][92] <= 18'h200ef;\
    linear1_weight_array[11][93] <= 18'h00121;\
    linear1_weight_array[11][94] <= 18'h000ba;\
    linear1_weight_array[11][95] <= 18'h00157;\
    linear1_weight_array[11][96] <= 18'h000e9;\
    linear1_weight_array[11][97] <= 18'h000aa;\
    linear1_weight_array[11][98] <= 18'h00041;\
    linear1_weight_array[11][99] <= 18'h000a3;\
    linear1_weight_array[11][100] <= 18'h0004c;\
    linear1_weight_array[11][101] <= 18'h200ea;\
    linear1_weight_array[11][102] <= 18'h2008b;\
    linear1_weight_array[11][103] <= 18'h2001c;\
    linear1_weight_array[11][104] <= 18'h00132;\
    linear1_weight_array[11][105] <= 18'h200ca;\
    linear1_weight_array[11][106] <= 18'h200fb;\
    linear1_weight_array[11][107] <= 18'h0000f;\
    linear1_weight_array[11][108] <= 18'h0002e;\
    linear1_weight_array[11][109] <= 18'h0007b;\
    linear1_weight_array[11][110] <= 18'h0002c;\
    linear1_weight_array[11][111] <= 18'h2006c;\
    linear1_weight_array[11][112] <= 18'h000c1;\
    linear1_weight_array[11][113] <= 18'h20084;\
    linear1_weight_array[11][114] <= 18'h20050;\
    linear1_weight_array[11][115] <= 18'h20092;\
    linear1_weight_array[11][116] <= 18'h00050;\
    linear1_weight_array[11][117] <= 18'h00064;\
    linear1_weight_array[11][118] <= 18'h0005a;\
    linear1_weight_array[11][119] <= 18'h0001f;\
    linear1_weight_array[11][120] <= 18'h00036;\
    linear1_weight_array[11][121] <= 18'h00022;\
    linear1_weight_array[11][122] <= 18'h0009d;\
    linear1_weight_array[11][123] <= 18'h00053;\
    linear1_weight_array[11][124] <= 18'h200b0;\
    linear1_weight_array[11][125] <= 18'h00229;\
    linear1_weight_array[11][126] <= 18'h000ad;\
    linear1_weight_array[11][127] <= 18'h0001a;\
    linear1_weight_array[11][128] <= 18'h2023a;\
    linear1_weight_array[11][129] <= 18'h202d9;\
    linear1_weight_array[11][130] <= 18'h0010a;\
    linear1_weight_array[11][131] <= 18'h00098;\
    linear1_weight_array[11][132] <= 18'h20059;\
    linear1_weight_array[11][133] <= 18'h20023;\
    linear1_weight_array[11][134] <= 18'h20148;\
    linear1_weight_array[11][135] <= 18'h200e6;\
    linear1_weight_array[11][136] <= 18'h00118;\
    linear1_weight_array[11][137] <= 18'h000a0;\
    linear1_weight_array[11][138] <= 18'h200fe;\
    linear1_weight_array[11][139] <= 18'h0004e;\
    linear1_weight_array[11][140] <= 18'h0007d;\
    linear1_weight_array[11][141] <= 18'h000dd;\
    linear1_weight_array[11][142] <= 18'h20023;\
    linear1_weight_array[11][143] <= 18'h20021;\
    linear1_weight_array[11][144] <= 18'h000d8;\
    linear1_weight_array[11][145] <= 18'h00055;\
    linear1_weight_array[11][146] <= 18'h00001;\
    linear1_weight_array[11][147] <= 18'h00019;\
    linear1_weight_array[11][148] <= 18'h0003c;\
    linear1_weight_array[11][149] <= 18'h20009;\
end

/*
`define LINEAR1_WEIGHT \
reg [0:17] linear1_weight_array [0:11][0:149];\
always@(posedge clk or negedge rst_n) begin\
    linear1_weight_array[0][0] <= 18'h00400;\
    linear1_weight_array[0][1] <= 18'h00600;\
    linear1_weight_array[0][2] <= 18'h20c00;\
    linear1_weight_array[0][3] <= 18'h00300;\
    linear1_weight_array[0][4] <= 18'h20080;\
    linear1_weight_array[0][5] <= 18'h00400;\
    linear1_weight_array[0][6] <= 18'h00600;\
    linear1_weight_array[0][7] <= 18'h20c00;\
    linear1_weight_array[0][8] <= 18'h00300;\
    linear1_weight_array[0][9] <= 18'h20080;\
    linear1_weight_array[0][10] <= 18'h00400;\
    linear1_weight_array[0][11] <= 18'h00600;\
    linear1_weight_array[0][12] <= 18'h20c00;\
    linear1_weight_array[0][13] <= 18'h00300;\
    linear1_weight_array[0][14] <= 18'h20080;\
    linear1_weight_array[0][15] <= 18'h00400;\
    linear1_weight_array[0][16] <= 18'h00600;\
    linear1_weight_array[0][17] <= 18'h20c00;\
    linear1_weight_array[0][18] <= 18'h00300;\
    linear1_weight_array[0][19] <= 18'h20080;\
    linear1_weight_array[0][20] <= 18'h00400;\
    linear1_weight_array[0][21] <= 18'h00600;\
    linear1_weight_array[0][22] <= 18'h20c00;\
    linear1_weight_array[0][23] <= 18'h00300;\
    linear1_weight_array[0][24] <= 18'h20080;\
    linear1_weight_array[0][25] <= 18'h00400;\
    linear1_weight_array[0][26] <= 18'h00600;\
    linear1_weight_array[0][27] <= 18'h20c00;\
    linear1_weight_array[0][28] <= 18'h00300;\
    linear1_weight_array[0][29] <= 18'h20080;\
    linear1_weight_array[0][30] <= 18'h00400;\
    linear1_weight_array[0][31] <= 18'h00600;\
    linear1_weight_array[0][32] <= 18'h20c00;\
    linear1_weight_array[0][33] <= 18'h00300;\
    linear1_weight_array[0][34] <= 18'h20080;\
    linear1_weight_array[0][35] <= 18'h00400;\
    linear1_weight_array[0][36] <= 18'h00600;\
    linear1_weight_array[0][37] <= 18'h20c00;\
    linear1_weight_array[0][38] <= 18'h00300;\
    linear1_weight_array[0][39] <= 18'h20080;\
    linear1_weight_array[0][40] <= 18'h00400;\
    linear1_weight_array[0][41] <= 18'h00600;\
    linear1_weight_array[0][42] <= 18'h20c00;\
    linear1_weight_array[0][43] <= 18'h00300;\
    linear1_weight_array[0][44] <= 18'h20080;\
    linear1_weight_array[0][45] <= 18'h00400;\
    linear1_weight_array[0][46] <= 18'h00600;\
    linear1_weight_array[0][47] <= 18'h20c00;\
    linear1_weight_array[0][48] <= 18'h00300;\
    linear1_weight_array[0][49] <= 18'h20080;\
    linear1_weight_array[0][50] <= 18'h00400;\
    linear1_weight_array[0][51] <= 18'h00600;\
    linear1_weight_array[0][52] <= 18'h20c00;\
    linear1_weight_array[0][53] <= 18'h00300;\
    linear1_weight_array[0][54] <= 18'h20080;\
    linear1_weight_array[0][55] <= 18'h00400;\
    linear1_weight_array[0][56] <= 18'h00600;\
    linear1_weight_array[0][57] <= 18'h20c00;\
    linear1_weight_array[0][58] <= 18'h00300;\
    linear1_weight_array[0][59] <= 18'h20080;\
    linear1_weight_array[0][60] <= 18'h00400;\
    linear1_weight_array[0][61] <= 18'h00600;\
    linear1_weight_array[0][62] <= 18'h20c00;\
    linear1_weight_array[0][63] <= 18'h00300;\
    linear1_weight_array[0][64] <= 18'h20080;\
    linear1_weight_array[0][65] <= 18'h00400;\
    linear1_weight_array[0][66] <= 18'h00600;\
    linear1_weight_array[0][67] <= 18'h20c00;\
    linear1_weight_array[0][68] <= 18'h00300;\
    linear1_weight_array[0][69] <= 18'h20080;\
    linear1_weight_array[0][70] <= 18'h00400;\
    linear1_weight_array[0][71] <= 18'h00600;\
    linear1_weight_array[0][72] <= 18'h20c00;\
    linear1_weight_array[0][73] <= 18'h00300;\
    linear1_weight_array[0][74] <= 18'h20080;\
    linear1_weight_array[0][75] <= 18'h00400;\
    linear1_weight_array[0][76] <= 18'h00600;\
    linear1_weight_array[0][77] <= 18'h20c00;\
    linear1_weight_array[0][78] <= 18'h00300;\
    linear1_weight_array[0][79] <= 18'h20080;\
    linear1_weight_array[0][80] <= 18'h00400;\
    linear1_weight_array[0][81] <= 18'h00600;\
    linear1_weight_array[0][82] <= 18'h20c00;\
    linear1_weight_array[0][83] <= 18'h00300;\
    linear1_weight_array[0][84] <= 18'h20080;\
    linear1_weight_array[0][85] <= 18'h00400;\
    linear1_weight_array[0][86] <= 18'h00600;\
    linear1_weight_array[0][87] <= 18'h20c00;\
    linear1_weight_array[0][88] <= 18'h00300;\
    linear1_weight_array[0][89] <= 18'h20080;\
    linear1_weight_array[0][90] <= 18'h00400;\
    linear1_weight_array[0][91] <= 18'h00600;\
    linear1_weight_array[0][92] <= 18'h20c00;\
    linear1_weight_array[0][93] <= 18'h00300;\
    linear1_weight_array[0][94] <= 18'h20080;\
    linear1_weight_array[0][95] <= 18'h00400;\
    linear1_weight_array[0][96] <= 18'h00600;\
    linear1_weight_array[0][97] <= 18'h20c00;\
    linear1_weight_array[0][98] <= 18'h00300;\
    linear1_weight_array[0][99] <= 18'h20080;\
    linear1_weight_array[0][100] <= 18'h00400;\
    linear1_weight_array[0][101] <= 18'h00600;\
    linear1_weight_array[0][102] <= 18'h20c00;\
    linear1_weight_array[0][103] <= 18'h00300;\
    linear1_weight_array[0][104] <= 18'h20080;\
    linear1_weight_array[0][105] <= 18'h00400;\
    linear1_weight_array[0][106] <= 18'h00600;\
    linear1_weight_array[0][107] <= 18'h20c00;\
    linear1_weight_array[0][108] <= 18'h00300;\
    linear1_weight_array[0][109] <= 18'h20080;\
    linear1_weight_array[0][110] <= 18'h00400;\
    linear1_weight_array[0][111] <= 18'h00600;\
    linear1_weight_array[0][112] <= 18'h20c00;\
    linear1_weight_array[0][113] <= 18'h00300;\
    linear1_weight_array[0][114] <= 18'h20080;\
    linear1_weight_array[0][115] <= 18'h00400;\
    linear1_weight_array[0][116] <= 18'h00600;\
    linear1_weight_array[0][117] <= 18'h20c00;\
    linear1_weight_array[0][118] <= 18'h00300;\
    linear1_weight_array[0][119] <= 18'h20080;\
    linear1_weight_array[0][120] <= 18'h00400;\
    linear1_weight_array[0][121] <= 18'h00600;\
    linear1_weight_array[0][122] <= 18'h20c00;\
    linear1_weight_array[0][123] <= 18'h00300;\
    linear1_weight_array[0][124] <= 18'h20080;\
    linear1_weight_array[0][125] <= 18'h00400;\
    linear1_weight_array[0][126] <= 18'h00600;\
    linear1_weight_array[0][127] <= 18'h20c00;\
    linear1_weight_array[0][128] <= 18'h00300;\
    linear1_weight_array[0][129] <= 18'h20080;\
    linear1_weight_array[0][130] <= 18'h00400;\
    linear1_weight_array[0][131] <= 18'h00600;\
    linear1_weight_array[0][132] <= 18'h20c00;\
    linear1_weight_array[0][133] <= 18'h00300;\
    linear1_weight_array[0][134] <= 18'h20080;\
    linear1_weight_array[0][135] <= 18'h00400;\
    linear1_weight_array[0][136] <= 18'h00600;\
    linear1_weight_array[0][137] <= 18'h20c00;\
    linear1_weight_array[0][138] <= 18'h00300;\
    linear1_weight_array[0][139] <= 18'h20080;\
    linear1_weight_array[0][140] <= 18'h00400;\
    linear1_weight_array[0][141] <= 18'h00600;\
    linear1_weight_array[0][142] <= 18'h20c00;\
    linear1_weight_array[0][143] <= 18'h00300;\
    linear1_weight_array[0][144] <= 18'h20080;\
    linear1_weight_array[0][145] <= 18'h00400;\
    linear1_weight_array[0][146] <= 18'h00600;\
    linear1_weight_array[0][147] <= 18'h20c00;\
    linear1_weight_array[0][148] <= 18'h00300;\
    linear1_weight_array[0][149] <= 18'h20080;\
    linear1_weight_array[1][0] <= 18'h00400;\
    linear1_weight_array[1][1] <= 18'h00600;\
    linear1_weight_array[1][2] <= 18'h20c00;\
    linear1_weight_array[1][3] <= 18'h00100;\
    linear1_weight_array[1][4] <= 18'h20080;\
    linear1_weight_array[1][5] <= 18'h00400;\
    linear1_weight_array[1][6] <= 18'h00600;\
    linear1_weight_array[1][7] <= 18'h20c00;\
    linear1_weight_array[1][8] <= 18'h00100;\
    linear1_weight_array[1][9] <= 18'h20080;\
    linear1_weight_array[1][10] <= 18'h00400;\
    linear1_weight_array[1][11] <= 18'h00600;\
    linear1_weight_array[1][12] <= 18'h20c00;\
    linear1_weight_array[1][13] <= 18'h00100;\
    linear1_weight_array[1][14] <= 18'h20080;\
    linear1_weight_array[1][15] <= 18'h00400;\
    linear1_weight_array[1][16] <= 18'h00600;\
    linear1_weight_array[1][17] <= 18'h20c00;\
    linear1_weight_array[1][18] <= 18'h00100;\
    linear1_weight_array[1][19] <= 18'h20080;\
    linear1_weight_array[1][20] <= 18'h00400;\
    linear1_weight_array[1][21] <= 18'h00600;\
    linear1_weight_array[1][22] <= 18'h20c00;\
    linear1_weight_array[1][23] <= 18'h00100;\
    linear1_weight_array[1][24] <= 18'h20080;\
    linear1_weight_array[1][25] <= 18'h00400;\
    linear1_weight_array[1][26] <= 18'h00600;\
    linear1_weight_array[1][27] <= 18'h20c00;\
    linear1_weight_array[1][28] <= 18'h00100;\
    linear1_weight_array[1][29] <= 18'h20080;\
    linear1_weight_array[1][30] <= 18'h00400;\
    linear1_weight_array[1][31] <= 18'h00600;\
    linear1_weight_array[1][32] <= 18'h20c00;\
    linear1_weight_array[1][33] <= 18'h00100;\
    linear1_weight_array[1][34] <= 18'h20080;\
    linear1_weight_array[1][35] <= 18'h00400;\
    linear1_weight_array[1][36] <= 18'h00600;\
    linear1_weight_array[1][37] <= 18'h20c00;\
    linear1_weight_array[1][38] <= 18'h00100;\
    linear1_weight_array[1][39] <= 18'h20080;\
    linear1_weight_array[1][40] <= 18'h00400;\
    linear1_weight_array[1][41] <= 18'h00600;\
    linear1_weight_array[1][42] <= 18'h20c00;\
    linear1_weight_array[1][43] <= 18'h00100;\
    linear1_weight_array[1][44] <= 18'h20080;\
    linear1_weight_array[1][45] <= 18'h00400;\
    linear1_weight_array[1][46] <= 18'h00600;\
    linear1_weight_array[1][47] <= 18'h20c00;\
    linear1_weight_array[1][48] <= 18'h00100;\
    linear1_weight_array[1][49] <= 18'h20080;\
    linear1_weight_array[1][50] <= 18'h00400;\
    linear1_weight_array[1][51] <= 18'h00600;\
    linear1_weight_array[1][52] <= 18'h20c00;\
    linear1_weight_array[1][53] <= 18'h00100;\
    linear1_weight_array[1][54] <= 18'h20080;\
    linear1_weight_array[1][55] <= 18'h00400;\
    linear1_weight_array[1][56] <= 18'h00600;\
    linear1_weight_array[1][57] <= 18'h20c00;\
    linear1_weight_array[1][58] <= 18'h00100;\
    linear1_weight_array[1][59] <= 18'h20080;\
    linear1_weight_array[1][60] <= 18'h00400;\
    linear1_weight_array[1][61] <= 18'h00600;\
    linear1_weight_array[1][62] <= 18'h20c00;\
    linear1_weight_array[1][63] <= 18'h00100;\
    linear1_weight_array[1][64] <= 18'h20080;\
    linear1_weight_array[1][65] <= 18'h00400;\
    linear1_weight_array[1][66] <= 18'h00600;\
    linear1_weight_array[1][67] <= 18'h20c00;\
    linear1_weight_array[1][68] <= 18'h00100;\
    linear1_weight_array[1][69] <= 18'h20080;\
    linear1_weight_array[1][70] <= 18'h00400;\
    linear1_weight_array[1][71] <= 18'h00600;\
    linear1_weight_array[1][72] <= 18'h20c00;\
    linear1_weight_array[1][73] <= 18'h00100;\
    linear1_weight_array[1][74] <= 18'h20080;\
    linear1_weight_array[1][75] <= 18'h00400;\
    linear1_weight_array[1][76] <= 18'h00600;\
    linear1_weight_array[1][77] <= 18'h20c00;\
    linear1_weight_array[1][78] <= 18'h00100;\
    linear1_weight_array[1][79] <= 18'h20080;\
    linear1_weight_array[1][80] <= 18'h00400;\
    linear1_weight_array[1][81] <= 18'h00600;\
    linear1_weight_array[1][82] <= 18'h20c00;\
    linear1_weight_array[1][83] <= 18'h00100;\
    linear1_weight_array[1][84] <= 18'h20080;\
    linear1_weight_array[1][85] <= 18'h00400;\
    linear1_weight_array[1][86] <= 18'h00600;\
    linear1_weight_array[1][87] <= 18'h20c00;\
    linear1_weight_array[1][88] <= 18'h00100;\
    linear1_weight_array[1][89] <= 18'h20080;\
    linear1_weight_array[1][90] <= 18'h00400;\
    linear1_weight_array[1][91] <= 18'h00600;\
    linear1_weight_array[1][92] <= 18'h20c00;\
    linear1_weight_array[1][93] <= 18'h00100;\
    linear1_weight_array[1][94] <= 18'h20080;\
    linear1_weight_array[1][95] <= 18'h00400;\
    linear1_weight_array[1][96] <= 18'h00600;\
    linear1_weight_array[1][97] <= 18'h20c00;\
    linear1_weight_array[1][98] <= 18'h00100;\
    linear1_weight_array[1][99] <= 18'h20080;\
    linear1_weight_array[1][100] <= 18'h00400;\
    linear1_weight_array[1][101] <= 18'h00600;\
    linear1_weight_array[1][102] <= 18'h20c00;\
    linear1_weight_array[1][103] <= 18'h00100;\
    linear1_weight_array[1][104] <= 18'h20080;\
    linear1_weight_array[1][105] <= 18'h00400;\
    linear1_weight_array[1][106] <= 18'h00600;\
    linear1_weight_array[1][107] <= 18'h20c00;\
    linear1_weight_array[1][108] <= 18'h00100;\
    linear1_weight_array[1][109] <= 18'h20080;\
    linear1_weight_array[1][110] <= 18'h00400;\
    linear1_weight_array[1][111] <= 18'h00600;\
    linear1_weight_array[1][112] <= 18'h20c00;\
    linear1_weight_array[1][113] <= 18'h00100;\
    linear1_weight_array[1][114] <= 18'h20080;\
    linear1_weight_array[1][115] <= 18'h00400;\
    linear1_weight_array[1][116] <= 18'h00600;\
    linear1_weight_array[1][117] <= 18'h20c00;\
    linear1_weight_array[1][118] <= 18'h00100;\
    linear1_weight_array[1][119] <= 18'h20080;\
    linear1_weight_array[1][120] <= 18'h00400;\
    linear1_weight_array[1][121] <= 18'h00600;\
    linear1_weight_array[1][122] <= 18'h20c00;\
    linear1_weight_array[1][123] <= 18'h00100;\
    linear1_weight_array[1][124] <= 18'h20080;\
    linear1_weight_array[1][125] <= 18'h00400;\
    linear1_weight_array[1][126] <= 18'h00600;\
    linear1_weight_array[1][127] <= 18'h20c00;\
    linear1_weight_array[1][128] <= 18'h00100;\
    linear1_weight_array[1][129] <= 18'h20080;\
    linear1_weight_array[1][130] <= 18'h00400;\
    linear1_weight_array[1][131] <= 18'h00600;\
    linear1_weight_array[1][132] <= 18'h20c00;\
    linear1_weight_array[1][133] <= 18'h00100;\
    linear1_weight_array[1][134] <= 18'h20080;\
    linear1_weight_array[1][135] <= 18'h00400;\
    linear1_weight_array[1][136] <= 18'h00600;\
    linear1_weight_array[1][137] <= 18'h20c00;\
    linear1_weight_array[1][138] <= 18'h00100;\
    linear1_weight_array[1][139] <= 18'h20080;\
    linear1_weight_array[1][140] <= 18'h00400;\
    linear1_weight_array[1][141] <= 18'h00600;\
    linear1_weight_array[1][142] <= 18'h20c00;\
    linear1_weight_array[1][143] <= 18'h00100;\
    linear1_weight_array[1][144] <= 18'h20080;\
    linear1_weight_array[1][145] <= 18'h00400;\
    linear1_weight_array[1][146] <= 18'h00600;\
    linear1_weight_array[1][147] <= 18'h20c00;\
    linear1_weight_array[1][148] <= 18'h00100;\
    linear1_weight_array[1][149] <= 18'h20080;\
    linear1_weight_array[2][0] <= 18'h00400;\
    linear1_weight_array[2][1] <= 18'h00600;\
    linear1_weight_array[2][2] <= 18'h20c00;\
    linear1_weight_array[2][3] <= 18'h00300;\
    linear1_weight_array[2][4] <= 18'h20080;\
    linear1_weight_array[2][5] <= 18'h00400;\
    linear1_weight_array[2][6] <= 18'h00600;\
    linear1_weight_array[2][7] <= 18'h20c00;\
    linear1_weight_array[2][8] <= 18'h00300;\
    linear1_weight_array[2][9] <= 18'h20080;\
    linear1_weight_array[2][10] <= 18'h00400;\
    linear1_weight_array[2][11] <= 18'h00600;\
    linear1_weight_array[2][12] <= 18'h20c00;\
    linear1_weight_array[2][13] <= 18'h00300;\
    linear1_weight_array[2][14] <= 18'h20080;\
    linear1_weight_array[2][15] <= 18'h00400;\
    linear1_weight_array[2][16] <= 18'h00600;\
    linear1_weight_array[2][17] <= 18'h20c00;\
    linear1_weight_array[2][18] <= 18'h00300;\
    linear1_weight_array[2][19] <= 18'h20080;\
    linear1_weight_array[2][20] <= 18'h00400;\
    linear1_weight_array[2][21] <= 18'h00600;\
    linear1_weight_array[2][22] <= 18'h20c00;\
    linear1_weight_array[2][23] <= 18'h00300;\
    linear1_weight_array[2][24] <= 18'h20080;\
    linear1_weight_array[2][25] <= 18'h00400;\
    linear1_weight_array[2][26] <= 18'h00600;\
    linear1_weight_array[2][27] <= 18'h20c00;\
    linear1_weight_array[2][28] <= 18'h00300;\
    linear1_weight_array[2][29] <= 18'h20080;\
    linear1_weight_array[2][30] <= 18'h00400;\
    linear1_weight_array[2][31] <= 18'h00600;\
    linear1_weight_array[2][32] <= 18'h20c00;\
    linear1_weight_array[2][33] <= 18'h00300;\
    linear1_weight_array[2][34] <= 18'h20080;\
    linear1_weight_array[2][35] <= 18'h00400;\
    linear1_weight_array[2][36] <= 18'h00600;\
    linear1_weight_array[2][37] <= 18'h20c00;\
    linear1_weight_array[2][38] <= 18'h00300;\
    linear1_weight_array[2][39] <= 18'h20080;\
    linear1_weight_array[2][40] <= 18'h00400;\
    linear1_weight_array[2][41] <= 18'h00600;\
    linear1_weight_array[2][42] <= 18'h20c00;\
    linear1_weight_array[2][43] <= 18'h00300;\
    linear1_weight_array[2][44] <= 18'h20080;\
    linear1_weight_array[2][45] <= 18'h00400;\
    linear1_weight_array[2][46] <= 18'h00600;\
    linear1_weight_array[2][47] <= 18'h20c00;\
    linear1_weight_array[2][48] <= 18'h00300;\
    linear1_weight_array[2][49] <= 18'h20080;\
    linear1_weight_array[2][50] <= 18'h00400;\
    linear1_weight_array[2][51] <= 18'h00600;\
    linear1_weight_array[2][52] <= 18'h20c00;\
    linear1_weight_array[2][53] <= 18'h00300;\
    linear1_weight_array[2][54] <= 18'h20080;\
    linear1_weight_array[2][55] <= 18'h00400;\
    linear1_weight_array[2][56] <= 18'h00600;\
    linear1_weight_array[2][57] <= 18'h20c00;\
    linear1_weight_array[2][58] <= 18'h00300;\
    linear1_weight_array[2][59] <= 18'h20080;\
    linear1_weight_array[2][60] <= 18'h00400;\
    linear1_weight_array[2][61] <= 18'h00600;\
    linear1_weight_array[2][62] <= 18'h20c00;\
    linear1_weight_array[2][63] <= 18'h00300;\
    linear1_weight_array[2][64] <= 18'h20080;\
    linear1_weight_array[2][65] <= 18'h00400;\
    linear1_weight_array[2][66] <= 18'h00600;\
    linear1_weight_array[2][67] <= 18'h20c00;\
    linear1_weight_array[2][68] <= 18'h00300;\
    linear1_weight_array[2][69] <= 18'h20080;\
    linear1_weight_array[2][70] <= 18'h00400;\
    linear1_weight_array[2][71] <= 18'h00600;\
    linear1_weight_array[2][72] <= 18'h20c00;\
    linear1_weight_array[2][73] <= 18'h00300;\
    linear1_weight_array[2][74] <= 18'h20080;\
    linear1_weight_array[2][75] <= 18'h00400;\
    linear1_weight_array[2][76] <= 18'h00600;\
    linear1_weight_array[2][77] <= 18'h20c00;\
    linear1_weight_array[2][78] <= 18'h00300;\
    linear1_weight_array[2][79] <= 18'h20080;\
    linear1_weight_array[2][80] <= 18'h00400;\
    linear1_weight_array[2][81] <= 18'h00600;\
    linear1_weight_array[2][82] <= 18'h20c00;\
    linear1_weight_array[2][83] <= 18'h00300;\
    linear1_weight_array[2][84] <= 18'h20080;\
    linear1_weight_array[2][85] <= 18'h00400;\
    linear1_weight_array[2][86] <= 18'h00600;\
    linear1_weight_array[2][87] <= 18'h20c00;\
    linear1_weight_array[2][88] <= 18'h00300;\
    linear1_weight_array[2][89] <= 18'h20080;\
    linear1_weight_array[2][90] <= 18'h00400;\
    linear1_weight_array[2][91] <= 18'h00600;\
    linear1_weight_array[2][92] <= 18'h20c00;\
    linear1_weight_array[2][93] <= 18'h00300;\
    linear1_weight_array[2][94] <= 18'h20080;\
    linear1_weight_array[2][95] <= 18'h00400;\
    linear1_weight_array[2][96] <= 18'h00600;\
    linear1_weight_array[2][97] <= 18'h20c00;\
    linear1_weight_array[2][98] <= 18'h00300;\
    linear1_weight_array[2][99] <= 18'h20080;\
    linear1_weight_array[2][100] <= 18'h00400;\
    linear1_weight_array[2][101] <= 18'h00600;\
    linear1_weight_array[2][102] <= 18'h20c00;\
    linear1_weight_array[2][103] <= 18'h00300;\
    linear1_weight_array[2][104] <= 18'h20080;\
    linear1_weight_array[2][105] <= 18'h00400;\
    linear1_weight_array[2][106] <= 18'h00600;\
    linear1_weight_array[2][107] <= 18'h20c00;\
    linear1_weight_array[2][108] <= 18'h00300;\
    linear1_weight_array[2][109] <= 18'h20080;\
    linear1_weight_array[2][110] <= 18'h00400;\
    linear1_weight_array[2][111] <= 18'h00600;\
    linear1_weight_array[2][112] <= 18'h20c00;\
    linear1_weight_array[2][113] <= 18'h00300;\
    linear1_weight_array[2][114] <= 18'h20080;\
    linear1_weight_array[2][115] <= 18'h00400;\
    linear1_weight_array[2][116] <= 18'h00600;\
    linear1_weight_array[2][117] <= 18'h20c00;\
    linear1_weight_array[2][118] <= 18'h00300;\
    linear1_weight_array[2][119] <= 18'h20080;\
    linear1_weight_array[2][120] <= 18'h00400;\
    linear1_weight_array[2][121] <= 18'h00600;\
    linear1_weight_array[2][122] <= 18'h20c00;\
    linear1_weight_array[2][123] <= 18'h00300;\
    linear1_weight_array[2][124] <= 18'h20080;\
    linear1_weight_array[2][125] <= 18'h00400;\
    linear1_weight_array[2][126] <= 18'h00600;\
    linear1_weight_array[2][127] <= 18'h20c00;\
    linear1_weight_array[2][128] <= 18'h00300;\
    linear1_weight_array[2][129] <= 18'h20080;\
    linear1_weight_array[2][130] <= 18'h00400;\
    linear1_weight_array[2][131] <= 18'h00600;\
    linear1_weight_array[2][132] <= 18'h20c00;\
    linear1_weight_array[2][133] <= 18'h00300;\
    linear1_weight_array[2][134] <= 18'h20080;\
    linear1_weight_array[2][135] <= 18'h00400;\
    linear1_weight_array[2][136] <= 18'h00600;\
    linear1_weight_array[2][137] <= 18'h20c00;\
    linear1_weight_array[2][138] <= 18'h00300;\
    linear1_weight_array[2][139] <= 18'h20080;\
    linear1_weight_array[2][140] <= 18'h00400;\
    linear1_weight_array[2][141] <= 18'h00600;\
    linear1_weight_array[2][142] <= 18'h20c00;\
    linear1_weight_array[2][143] <= 18'h00300;\
    linear1_weight_array[2][144] <= 18'h20080;\
    linear1_weight_array[2][145] <= 18'h00400;\
    linear1_weight_array[2][146] <= 18'h00600;\
    linear1_weight_array[2][147] <= 18'h20c00;\
    linear1_weight_array[2][148] <= 18'h00300;\
    linear1_weight_array[2][149] <= 18'h20080;\
    linear1_weight_array[3][0] <= 18'h00400;\
    linear1_weight_array[3][1] <= 18'h00600;\
    linear1_weight_array[3][2] <= 18'h20c00;\
    linear1_weight_array[3][3] <= 18'h00100;\
    linear1_weight_array[3][4] <= 18'h20080;\
    linear1_weight_array[3][5] <= 18'h00400;\
    linear1_weight_array[3][6] <= 18'h00600;\
    linear1_weight_array[3][7] <= 18'h20c00;\
    linear1_weight_array[3][8] <= 18'h00100;\
    linear1_weight_array[3][9] <= 18'h20080;\
    linear1_weight_array[3][10] <= 18'h00400;\
    linear1_weight_array[3][11] <= 18'h00600;\
    linear1_weight_array[3][12] <= 18'h20c00;\
    linear1_weight_array[3][13] <= 18'h00100;\
    linear1_weight_array[3][14] <= 18'h20080;\
    linear1_weight_array[3][15] <= 18'h00400;\
    linear1_weight_array[3][16] <= 18'h00600;\
    linear1_weight_array[3][17] <= 18'h20c00;\
    linear1_weight_array[3][18] <= 18'h00100;\
    linear1_weight_array[3][19] <= 18'h20080;\
    linear1_weight_array[3][20] <= 18'h00400;\
    linear1_weight_array[3][21] <= 18'h00600;\
    linear1_weight_array[3][22] <= 18'h20c00;\
    linear1_weight_array[3][23] <= 18'h00100;\
    linear1_weight_array[3][24] <= 18'h20080;\
    linear1_weight_array[3][25] <= 18'h00400;\
    linear1_weight_array[3][26] <= 18'h00600;\
    linear1_weight_array[3][27] <= 18'h20c00;\
    linear1_weight_array[3][28] <= 18'h00100;\
    linear1_weight_array[3][29] <= 18'h20080;\
    linear1_weight_array[3][30] <= 18'h00400;\
    linear1_weight_array[3][31] <= 18'h00600;\
    linear1_weight_array[3][32] <= 18'h20c00;\
    linear1_weight_array[3][33] <= 18'h00100;\
    linear1_weight_array[3][34] <= 18'h20080;\
    linear1_weight_array[3][35] <= 18'h00400;\
    linear1_weight_array[3][36] <= 18'h00600;\
    linear1_weight_array[3][37] <= 18'h20c00;\
    linear1_weight_array[3][38] <= 18'h00100;\
    linear1_weight_array[3][39] <= 18'h20080;\
    linear1_weight_array[3][40] <= 18'h00400;\
    linear1_weight_array[3][41] <= 18'h00600;\
    linear1_weight_array[3][42] <= 18'h20c00;\
    linear1_weight_array[3][43] <= 18'h00100;\
    linear1_weight_array[3][44] <= 18'h20080;\
    linear1_weight_array[3][45] <= 18'h00400;\
    linear1_weight_array[3][46] <= 18'h00600;\
    linear1_weight_array[3][47] <= 18'h20c00;\
    linear1_weight_array[3][48] <= 18'h00100;\
    linear1_weight_array[3][49] <= 18'h20080;\
    linear1_weight_array[3][50] <= 18'h00400;\
    linear1_weight_array[3][51] <= 18'h00600;\
    linear1_weight_array[3][52] <= 18'h20c00;\
    linear1_weight_array[3][53] <= 18'h00100;\
    linear1_weight_array[3][54] <= 18'h20080;\
    linear1_weight_array[3][55] <= 18'h00400;\
    linear1_weight_array[3][56] <= 18'h00600;\
    linear1_weight_array[3][57] <= 18'h20c00;\
    linear1_weight_array[3][58] <= 18'h00100;\
    linear1_weight_array[3][59] <= 18'h20080;\
    linear1_weight_array[3][60] <= 18'h00400;\
    linear1_weight_array[3][61] <= 18'h00600;\
    linear1_weight_array[3][62] <= 18'h20c00;\
    linear1_weight_array[3][63] <= 18'h00100;\
    linear1_weight_array[3][64] <= 18'h20080;\
    linear1_weight_array[3][65] <= 18'h00400;\
    linear1_weight_array[3][66] <= 18'h00600;\
    linear1_weight_array[3][67] <= 18'h20c00;\
    linear1_weight_array[3][68] <= 18'h00100;\
    linear1_weight_array[3][69] <= 18'h20080;\
    linear1_weight_array[3][70] <= 18'h00400;\
    linear1_weight_array[3][71] <= 18'h00600;\
    linear1_weight_array[3][72] <= 18'h20c00;\
    linear1_weight_array[3][73] <= 18'h00100;\
    linear1_weight_array[3][74] <= 18'h20080;\
    linear1_weight_array[3][75] <= 18'h00400;\
    linear1_weight_array[3][76] <= 18'h00600;\
    linear1_weight_array[3][77] <= 18'h20c00;\
    linear1_weight_array[3][78] <= 18'h00100;\
    linear1_weight_array[3][79] <= 18'h20080;\
    linear1_weight_array[3][80] <= 18'h00400;\
    linear1_weight_array[3][81] <= 18'h00600;\
    linear1_weight_array[3][82] <= 18'h20c00;\
    linear1_weight_array[3][83] <= 18'h00100;\
    linear1_weight_array[3][84] <= 18'h20080;\
    linear1_weight_array[3][85] <= 18'h00400;\
    linear1_weight_array[3][86] <= 18'h00600;\
    linear1_weight_array[3][87] <= 18'h20c00;\
    linear1_weight_array[3][88] <= 18'h00100;\
    linear1_weight_array[3][89] <= 18'h20080;\
    linear1_weight_array[3][90] <= 18'h00400;\
    linear1_weight_array[3][91] <= 18'h00600;\
    linear1_weight_array[3][92] <= 18'h20c00;\
    linear1_weight_array[3][93] <= 18'h00100;\
    linear1_weight_array[3][94] <= 18'h20080;\
    linear1_weight_array[3][95] <= 18'h00400;\
    linear1_weight_array[3][96] <= 18'h00600;\
    linear1_weight_array[3][97] <= 18'h20c00;\
    linear1_weight_array[3][98] <= 18'h00100;\
    linear1_weight_array[3][99] <= 18'h20080;\
    linear1_weight_array[3][100] <= 18'h00400;\
    linear1_weight_array[3][101] <= 18'h00600;\
    linear1_weight_array[3][102] <= 18'h20c00;\
    linear1_weight_array[3][103] <= 18'h00100;\
    linear1_weight_array[3][104] <= 18'h20080;\
    linear1_weight_array[3][105] <= 18'h00400;\
    linear1_weight_array[3][106] <= 18'h00600;\
    linear1_weight_array[3][107] <= 18'h20c00;\
    linear1_weight_array[3][108] <= 18'h00100;\
    linear1_weight_array[3][109] <= 18'h20080;\
    linear1_weight_array[3][110] <= 18'h00400;\
    linear1_weight_array[3][111] <= 18'h00600;\
    linear1_weight_array[3][112] <= 18'h20c00;\
    linear1_weight_array[3][113] <= 18'h00100;\
    linear1_weight_array[3][114] <= 18'h20080;\
    linear1_weight_array[3][115] <= 18'h00400;\
    linear1_weight_array[3][116] <= 18'h00600;\
    linear1_weight_array[3][117] <= 18'h20c00;\
    linear1_weight_array[3][118] <= 18'h00100;\
    linear1_weight_array[3][119] <= 18'h20080;\
    linear1_weight_array[3][120] <= 18'h00400;\
    linear1_weight_array[3][121] <= 18'h00600;\
    linear1_weight_array[3][122] <= 18'h20c00;\
    linear1_weight_array[3][123] <= 18'h00100;\
    linear1_weight_array[3][124] <= 18'h20080;\
    linear1_weight_array[3][125] <= 18'h00400;\
    linear1_weight_array[3][126] <= 18'h00600;\
    linear1_weight_array[3][127] <= 18'h20c00;\
    linear1_weight_array[3][128] <= 18'h00100;\
    linear1_weight_array[3][129] <= 18'h20080;\
    linear1_weight_array[3][130] <= 18'h00400;\
    linear1_weight_array[3][131] <= 18'h00600;\
    linear1_weight_array[3][132] <= 18'h20c00;\
    linear1_weight_array[3][133] <= 18'h00100;\
    linear1_weight_array[3][134] <= 18'h20080;\
    linear1_weight_array[3][135] <= 18'h00400;\
    linear1_weight_array[3][136] <= 18'h00600;\
    linear1_weight_array[3][137] <= 18'h20c00;\
    linear1_weight_array[3][138] <= 18'h00100;\
    linear1_weight_array[3][139] <= 18'h20080;\
    linear1_weight_array[3][140] <= 18'h00400;\
    linear1_weight_array[3][141] <= 18'h00600;\
    linear1_weight_array[3][142] <= 18'h20c00;\
    linear1_weight_array[3][143] <= 18'h00100;\
    linear1_weight_array[3][144] <= 18'h20080;\
    linear1_weight_array[3][145] <= 18'h00400;\
    linear1_weight_array[3][146] <= 18'h00600;\
    linear1_weight_array[3][147] <= 18'h20c00;\
    linear1_weight_array[3][148] <= 18'h00100;\
    linear1_weight_array[3][149] <= 18'h20080;\
    linear1_weight_array[4][0] <= 18'h00400;\
    linear1_weight_array[4][1] <= 18'h00600;\
    linear1_weight_array[4][2] <= 18'h20c00;\
    linear1_weight_array[4][3] <= 18'h00300;\
    linear1_weight_array[4][4] <= 18'h20080;\
    linear1_weight_array[4][5] <= 18'h00400;\
    linear1_weight_array[4][6] <= 18'h00600;\
    linear1_weight_array[4][7] <= 18'h20c00;\
    linear1_weight_array[4][8] <= 18'h00300;\
    linear1_weight_array[4][9] <= 18'h20080;\
    linear1_weight_array[4][10] <= 18'h00400;\
    linear1_weight_array[4][11] <= 18'h00600;\
    linear1_weight_array[4][12] <= 18'h20c00;\
    linear1_weight_array[4][13] <= 18'h00300;\
    linear1_weight_array[4][14] <= 18'h20080;\
    linear1_weight_array[4][15] <= 18'h00400;\
    linear1_weight_array[4][16] <= 18'h00600;\
    linear1_weight_array[4][17] <= 18'h20c00;\
    linear1_weight_array[4][18] <= 18'h00300;\
    linear1_weight_array[4][19] <= 18'h20080;\
    linear1_weight_array[4][20] <= 18'h00400;\
    linear1_weight_array[4][21] <= 18'h00600;\
    linear1_weight_array[4][22] <= 18'h20c00;\
    linear1_weight_array[4][23] <= 18'h00300;\
    linear1_weight_array[4][24] <= 18'h20080;\
    linear1_weight_array[4][25] <= 18'h00400;\
    linear1_weight_array[4][26] <= 18'h00600;\
    linear1_weight_array[4][27] <= 18'h20c00;\
    linear1_weight_array[4][28] <= 18'h00300;\
    linear1_weight_array[4][29] <= 18'h20080;\
    linear1_weight_array[4][30] <= 18'h00400;\
    linear1_weight_array[4][31] <= 18'h00600;\
    linear1_weight_array[4][32] <= 18'h20c00;\
    linear1_weight_array[4][33] <= 18'h00300;\
    linear1_weight_array[4][34] <= 18'h20080;\
    linear1_weight_array[4][35] <= 18'h00400;\
    linear1_weight_array[4][36] <= 18'h00600;\
    linear1_weight_array[4][37] <= 18'h20c00;\
    linear1_weight_array[4][38] <= 18'h00300;\
    linear1_weight_array[4][39] <= 18'h20080;\
    linear1_weight_array[4][40] <= 18'h00400;\
    linear1_weight_array[4][41] <= 18'h00600;\
    linear1_weight_array[4][42] <= 18'h20c00;\
    linear1_weight_array[4][43] <= 18'h00300;\
    linear1_weight_array[4][44] <= 18'h20080;\
    linear1_weight_array[4][45] <= 18'h00400;\
    linear1_weight_array[4][46] <= 18'h00600;\
    linear1_weight_array[4][47] <= 18'h20c00;\
    linear1_weight_array[4][48] <= 18'h00300;\
    linear1_weight_array[4][49] <= 18'h20080;\
    linear1_weight_array[4][50] <= 18'h00400;\
    linear1_weight_array[4][51] <= 18'h00600;\
    linear1_weight_array[4][52] <= 18'h20c00;\
    linear1_weight_array[4][53] <= 18'h00300;\
    linear1_weight_array[4][54] <= 18'h20080;\
    linear1_weight_array[4][55] <= 18'h00400;\
    linear1_weight_array[4][56] <= 18'h00600;\
    linear1_weight_array[4][57] <= 18'h20c00;\
    linear1_weight_array[4][58] <= 18'h00300;\
    linear1_weight_array[4][59] <= 18'h20080;\
    linear1_weight_array[4][60] <= 18'h00400;\
    linear1_weight_array[4][61] <= 18'h00600;\
    linear1_weight_array[4][62] <= 18'h20c00;\
    linear1_weight_array[4][63] <= 18'h00300;\
    linear1_weight_array[4][64] <= 18'h20080;\
    linear1_weight_array[4][65] <= 18'h00400;\
    linear1_weight_array[4][66] <= 18'h00600;\
    linear1_weight_array[4][67] <= 18'h20c00;\
    linear1_weight_array[4][68] <= 18'h00300;\
    linear1_weight_array[4][69] <= 18'h20080;\
    linear1_weight_array[4][70] <= 18'h00400;\
    linear1_weight_array[4][71] <= 18'h00600;\
    linear1_weight_array[4][72] <= 18'h20c00;\
    linear1_weight_array[4][73] <= 18'h00300;\
    linear1_weight_array[4][74] <= 18'h20080;\
    linear1_weight_array[4][75] <= 18'h00400;\
    linear1_weight_array[4][76] <= 18'h00600;\
    linear1_weight_array[4][77] <= 18'h20c00;\
    linear1_weight_array[4][78] <= 18'h00300;\
    linear1_weight_array[4][79] <= 18'h20080;\
    linear1_weight_array[4][80] <= 18'h00400;\
    linear1_weight_array[4][81] <= 18'h00600;\
    linear1_weight_array[4][82] <= 18'h20c00;\
    linear1_weight_array[4][83] <= 18'h00300;\
    linear1_weight_array[4][84] <= 18'h20080;\
    linear1_weight_array[4][85] <= 18'h00400;\
    linear1_weight_array[4][86] <= 18'h00600;\
    linear1_weight_array[4][87] <= 18'h20c00;\
    linear1_weight_array[4][88] <= 18'h00300;\
    linear1_weight_array[4][89] <= 18'h20080;\
    linear1_weight_array[4][90] <= 18'h00400;\
    linear1_weight_array[4][91] <= 18'h00600;\
    linear1_weight_array[4][92] <= 18'h20c00;\
    linear1_weight_array[4][93] <= 18'h00300;\
    linear1_weight_array[4][94] <= 18'h20080;\
    linear1_weight_array[4][95] <= 18'h00400;\
    linear1_weight_array[4][96] <= 18'h00600;\
    linear1_weight_array[4][97] <= 18'h20c00;\
    linear1_weight_array[4][98] <= 18'h00300;\
    linear1_weight_array[4][99] <= 18'h20080;\
    linear1_weight_array[4][100] <= 18'h00400;\
    linear1_weight_array[4][101] <= 18'h00600;\
    linear1_weight_array[4][102] <= 18'h20c00;\
    linear1_weight_array[4][103] <= 18'h00300;\
    linear1_weight_array[4][104] <= 18'h20080;\
    linear1_weight_array[4][105] <= 18'h00400;\
    linear1_weight_array[4][106] <= 18'h00600;\
    linear1_weight_array[4][107] <= 18'h20c00;\
    linear1_weight_array[4][108] <= 18'h00300;\
    linear1_weight_array[4][109] <= 18'h20080;\
    linear1_weight_array[4][110] <= 18'h00400;\
    linear1_weight_array[4][111] <= 18'h00600;\
    linear1_weight_array[4][112] <= 18'h20c00;\
    linear1_weight_array[4][113] <= 18'h00300;\
    linear1_weight_array[4][114] <= 18'h20080;\
    linear1_weight_array[4][115] <= 18'h00400;\
    linear1_weight_array[4][116] <= 18'h00600;\
    linear1_weight_array[4][117] <= 18'h20c00;\
    linear1_weight_array[4][118] <= 18'h00300;\
    linear1_weight_array[4][119] <= 18'h20080;\
    linear1_weight_array[4][120] <= 18'h00400;\
    linear1_weight_array[4][121] <= 18'h00600;\
    linear1_weight_array[4][122] <= 18'h20c00;\
    linear1_weight_array[4][123] <= 18'h00300;\
    linear1_weight_array[4][124] <= 18'h20080;\
    linear1_weight_array[4][125] <= 18'h00400;\
    linear1_weight_array[4][126] <= 18'h00600;\
    linear1_weight_array[4][127] <= 18'h20c00;\
    linear1_weight_array[4][128] <= 18'h00300;\
    linear1_weight_array[4][129] <= 18'h20080;\
    linear1_weight_array[4][130] <= 18'h00400;\
    linear1_weight_array[4][131] <= 18'h00600;\
    linear1_weight_array[4][132] <= 18'h20c00;\
    linear1_weight_array[4][133] <= 18'h00300;\
    linear1_weight_array[4][134] <= 18'h20080;\
    linear1_weight_array[4][135] <= 18'h00400;\
    linear1_weight_array[4][136] <= 18'h00600;\
    linear1_weight_array[4][137] <= 18'h20c00;\
    linear1_weight_array[4][138] <= 18'h00300;\
    linear1_weight_array[4][139] <= 18'h20080;\
    linear1_weight_array[4][140] <= 18'h00400;\
    linear1_weight_array[4][141] <= 18'h00600;\
    linear1_weight_array[4][142] <= 18'h20c00;\
    linear1_weight_array[4][143] <= 18'h00300;\
    linear1_weight_array[4][144] <= 18'h20080;\
    linear1_weight_array[4][145] <= 18'h00400;\
    linear1_weight_array[4][146] <= 18'h00600;\
    linear1_weight_array[4][147] <= 18'h20c00;\
    linear1_weight_array[4][148] <= 18'h00300;\
    linear1_weight_array[4][149] <= 18'h20080;\
    linear1_weight_array[5][0] <= 18'h00400;\
    linear1_weight_array[5][1] <= 18'h00600;\
    linear1_weight_array[5][2] <= 18'h20c00;\
    linear1_weight_array[5][3] <= 18'h00100;\
    linear1_weight_array[5][4] <= 18'h20080;\
    linear1_weight_array[5][5] <= 18'h00400;\
    linear1_weight_array[5][6] <= 18'h00600;\
    linear1_weight_array[5][7] <= 18'h20c00;\
    linear1_weight_array[5][8] <= 18'h00100;\
    linear1_weight_array[5][9] <= 18'h20080;\
    linear1_weight_array[5][10] <= 18'h00400;\
    linear1_weight_array[5][11] <= 18'h00600;\
    linear1_weight_array[5][12] <= 18'h20c00;\
    linear1_weight_array[5][13] <= 18'h00100;\
    linear1_weight_array[5][14] <= 18'h20080;\
    linear1_weight_array[5][15] <= 18'h00400;\
    linear1_weight_array[5][16] <= 18'h00600;\
    linear1_weight_array[5][17] <= 18'h20c00;\
    linear1_weight_array[5][18] <= 18'h00100;\
    linear1_weight_array[5][19] <= 18'h20080;\
    linear1_weight_array[5][20] <= 18'h00400;\
    linear1_weight_array[5][21] <= 18'h00600;\
    linear1_weight_array[5][22] <= 18'h20c00;\
    linear1_weight_array[5][23] <= 18'h00100;\
    linear1_weight_array[5][24] <= 18'h20080;\
    linear1_weight_array[5][25] <= 18'h00400;\
    linear1_weight_array[5][26] <= 18'h00600;\
    linear1_weight_array[5][27] <= 18'h20c00;\
    linear1_weight_array[5][28] <= 18'h00100;\
    linear1_weight_array[5][29] <= 18'h20080;\
    linear1_weight_array[5][30] <= 18'h00400;\
    linear1_weight_array[5][31] <= 18'h00600;\
    linear1_weight_array[5][32] <= 18'h20c00;\
    linear1_weight_array[5][33] <= 18'h00100;\
    linear1_weight_array[5][34] <= 18'h20080;\
    linear1_weight_array[5][35] <= 18'h00400;\
    linear1_weight_array[5][36] <= 18'h00600;\
    linear1_weight_array[5][37] <= 18'h20c00;\
    linear1_weight_array[5][38] <= 18'h00100;\
    linear1_weight_array[5][39] <= 18'h20080;\
    linear1_weight_array[5][40] <= 18'h00400;\
    linear1_weight_array[5][41] <= 18'h00600;\
    linear1_weight_array[5][42] <= 18'h20c00;\
    linear1_weight_array[5][43] <= 18'h00100;\
    linear1_weight_array[5][44] <= 18'h20080;\
    linear1_weight_array[5][45] <= 18'h00400;\
    linear1_weight_array[5][46] <= 18'h00600;\
    linear1_weight_array[5][47] <= 18'h20c00;\
    linear1_weight_array[5][48] <= 18'h00100;\
    linear1_weight_array[5][49] <= 18'h20080;\
    linear1_weight_array[5][50] <= 18'h00400;\
    linear1_weight_array[5][51] <= 18'h00600;\
    linear1_weight_array[5][52] <= 18'h20c00;\
    linear1_weight_array[5][53] <= 18'h00100;\
    linear1_weight_array[5][54] <= 18'h20080;\
    linear1_weight_array[5][55] <= 18'h00400;\
    linear1_weight_array[5][56] <= 18'h00600;\
    linear1_weight_array[5][57] <= 18'h20c00;\
    linear1_weight_array[5][58] <= 18'h00100;\
    linear1_weight_array[5][59] <= 18'h20080;\
    linear1_weight_array[5][60] <= 18'h00400;\
    linear1_weight_array[5][61] <= 18'h00600;\
    linear1_weight_array[5][62] <= 18'h20c00;\
    linear1_weight_array[5][63] <= 18'h00100;\
    linear1_weight_array[5][64] <= 18'h20080;\
    linear1_weight_array[5][65] <= 18'h00400;\
    linear1_weight_array[5][66] <= 18'h00600;\
    linear1_weight_array[5][67] <= 18'h20c00;\
    linear1_weight_array[5][68] <= 18'h00100;\
    linear1_weight_array[5][69] <= 18'h20080;\
    linear1_weight_array[5][70] <= 18'h00400;\
    linear1_weight_array[5][71] <= 18'h00600;\
    linear1_weight_array[5][72] <= 18'h20c00;\
    linear1_weight_array[5][73] <= 18'h00100;\
    linear1_weight_array[5][74] <= 18'h20080;\
    linear1_weight_array[5][75] <= 18'h00400;\
    linear1_weight_array[5][76] <= 18'h00600;\
    linear1_weight_array[5][77] <= 18'h20c00;\
    linear1_weight_array[5][78] <= 18'h00100;\
    linear1_weight_array[5][79] <= 18'h20080;\
    linear1_weight_array[5][80] <= 18'h00400;\
    linear1_weight_array[5][81] <= 18'h00600;\
    linear1_weight_array[5][82] <= 18'h20c00;\
    linear1_weight_array[5][83] <= 18'h00100;\
    linear1_weight_array[5][84] <= 18'h20080;\
    linear1_weight_array[5][85] <= 18'h00400;\
    linear1_weight_array[5][86] <= 18'h00600;\
    linear1_weight_array[5][87] <= 18'h20c00;\
    linear1_weight_array[5][88] <= 18'h00100;\
    linear1_weight_array[5][89] <= 18'h20080;\
    linear1_weight_array[5][90] <= 18'h00400;\
    linear1_weight_array[5][91] <= 18'h00600;\
    linear1_weight_array[5][92] <= 18'h20c00;\
    linear1_weight_array[5][93] <= 18'h00100;\
    linear1_weight_array[5][94] <= 18'h20080;\
    linear1_weight_array[5][95] <= 18'h00400;\
    linear1_weight_array[5][96] <= 18'h00600;\
    linear1_weight_array[5][97] <= 18'h20c00;\
    linear1_weight_array[5][98] <= 18'h00100;\
    linear1_weight_array[5][99] <= 18'h20080;\
    linear1_weight_array[5][100] <= 18'h00400;\
    linear1_weight_array[5][101] <= 18'h00600;\
    linear1_weight_array[5][102] <= 18'h20c00;\
    linear1_weight_array[5][103] <= 18'h00100;\
    linear1_weight_array[5][104] <= 18'h20080;\
    linear1_weight_array[5][105] <= 18'h00400;\
    linear1_weight_array[5][106] <= 18'h00600;\
    linear1_weight_array[5][107] <= 18'h20c00;\
    linear1_weight_array[5][108] <= 18'h00100;\
    linear1_weight_array[5][109] <= 18'h20080;\
    linear1_weight_array[5][110] <= 18'h00400;\
    linear1_weight_array[5][111] <= 18'h00600;\
    linear1_weight_array[5][112] <= 18'h20c00;\
    linear1_weight_array[5][113] <= 18'h00100;\
    linear1_weight_array[5][114] <= 18'h20080;\
    linear1_weight_array[5][115] <= 18'h00400;\
    linear1_weight_array[5][116] <= 18'h00600;\
    linear1_weight_array[5][117] <= 18'h20c00;\
    linear1_weight_array[5][118] <= 18'h00100;\
    linear1_weight_array[5][119] <= 18'h20080;\
    linear1_weight_array[5][120] <= 18'h00400;\
    linear1_weight_array[5][121] <= 18'h00600;\
    linear1_weight_array[5][122] <= 18'h20c00;\
    linear1_weight_array[5][123] <= 18'h00100;\
    linear1_weight_array[5][124] <= 18'h20080;\
    linear1_weight_array[5][125] <= 18'h00400;\
    linear1_weight_array[5][126] <= 18'h00600;\
    linear1_weight_array[5][127] <= 18'h20c00;\
    linear1_weight_array[5][128] <= 18'h00100;\
    linear1_weight_array[5][129] <= 18'h20080;\
    linear1_weight_array[5][130] <= 18'h00400;\
    linear1_weight_array[5][131] <= 18'h00600;\
    linear1_weight_array[5][132] <= 18'h20c00;\
    linear1_weight_array[5][133] <= 18'h00100;\
    linear1_weight_array[5][134] <= 18'h20080;\
    linear1_weight_array[5][135] <= 18'h00400;\
    linear1_weight_array[5][136] <= 18'h00600;\
    linear1_weight_array[5][137] <= 18'h20c00;\
    linear1_weight_array[5][138] <= 18'h00100;\
    linear1_weight_array[5][139] <= 18'h20080;\
    linear1_weight_array[5][140] <= 18'h00400;\
    linear1_weight_array[5][141] <= 18'h00600;\
    linear1_weight_array[5][142] <= 18'h20c00;\
    linear1_weight_array[5][143] <= 18'h00100;\
    linear1_weight_array[5][144] <= 18'h20080;\
    linear1_weight_array[5][145] <= 18'h00400;\
    linear1_weight_array[5][146] <= 18'h00600;\
    linear1_weight_array[5][147] <= 18'h20c00;\
    linear1_weight_array[5][148] <= 18'h00100;\
    linear1_weight_array[5][149] <= 18'h20080;\
    linear1_weight_array[6][0] <= 18'h00400;\
    linear1_weight_array[6][1] <= 18'h00600;\
    linear1_weight_array[6][2] <= 18'h20c00;\
    linear1_weight_array[6][3] <= 18'h00300;\
    linear1_weight_array[6][4] <= 18'h20080;\
    linear1_weight_array[6][5] <= 18'h00400;\
    linear1_weight_array[6][6] <= 18'h00600;\
    linear1_weight_array[6][7] <= 18'h20c00;\
    linear1_weight_array[6][8] <= 18'h00300;\
    linear1_weight_array[6][9] <= 18'h20080;\
    linear1_weight_array[6][10] <= 18'h00400;\
    linear1_weight_array[6][11] <= 18'h00600;\
    linear1_weight_array[6][12] <= 18'h20c00;\
    linear1_weight_array[6][13] <= 18'h00300;\
    linear1_weight_array[6][14] <= 18'h20080;\
    linear1_weight_array[6][15] <= 18'h00400;\
    linear1_weight_array[6][16] <= 18'h00600;\
    linear1_weight_array[6][17] <= 18'h20c00;\
    linear1_weight_array[6][18] <= 18'h00300;\
    linear1_weight_array[6][19] <= 18'h20080;\
    linear1_weight_array[6][20] <= 18'h00400;\
    linear1_weight_array[6][21] <= 18'h00600;\
    linear1_weight_array[6][22] <= 18'h20c00;\
    linear1_weight_array[6][23] <= 18'h00300;\
    linear1_weight_array[6][24] <= 18'h20080;\
    linear1_weight_array[6][25] <= 18'h00400;\
    linear1_weight_array[6][26] <= 18'h00600;\
    linear1_weight_array[6][27] <= 18'h20c00;\
    linear1_weight_array[6][28] <= 18'h00300;\
    linear1_weight_array[6][29] <= 18'h20080;\
    linear1_weight_array[6][30] <= 18'h00400;\
    linear1_weight_array[6][31] <= 18'h00600;\
    linear1_weight_array[6][32] <= 18'h20c00;\
    linear1_weight_array[6][33] <= 18'h00300;\
    linear1_weight_array[6][34] <= 18'h20080;\
    linear1_weight_array[6][35] <= 18'h00400;\
    linear1_weight_array[6][36] <= 18'h00600;\
    linear1_weight_array[6][37] <= 18'h20c00;\
    linear1_weight_array[6][38] <= 18'h00300;\
    linear1_weight_array[6][39] <= 18'h20080;\
    linear1_weight_array[6][40] <= 18'h00400;\
    linear1_weight_array[6][41] <= 18'h00600;\
    linear1_weight_array[6][42] <= 18'h20c00;\
    linear1_weight_array[6][43] <= 18'h00300;\
    linear1_weight_array[6][44] <= 18'h20080;\
    linear1_weight_array[6][45] <= 18'h00400;\
    linear1_weight_array[6][46] <= 18'h00600;\
    linear1_weight_array[6][47] <= 18'h20c00;\
    linear1_weight_array[6][48] <= 18'h00300;\
    linear1_weight_array[6][49] <= 18'h20080;\
    linear1_weight_array[6][50] <= 18'h00400;\
    linear1_weight_array[6][51] <= 18'h00600;\
    linear1_weight_array[6][52] <= 18'h20c00;\
    linear1_weight_array[6][53] <= 18'h00300;\
    linear1_weight_array[6][54] <= 18'h20080;\
    linear1_weight_array[6][55] <= 18'h00400;\
    linear1_weight_array[6][56] <= 18'h00600;\
    linear1_weight_array[6][57] <= 18'h20c00;\
    linear1_weight_array[6][58] <= 18'h00300;\
    linear1_weight_array[6][59] <= 18'h20080;\
    linear1_weight_array[6][60] <= 18'h00400;\
    linear1_weight_array[6][61] <= 18'h00600;\
    linear1_weight_array[6][62] <= 18'h20c00;\
    linear1_weight_array[6][63] <= 18'h00300;\
    linear1_weight_array[6][64] <= 18'h20080;\
    linear1_weight_array[6][65] <= 18'h00400;\
    linear1_weight_array[6][66] <= 18'h00600;\
    linear1_weight_array[6][67] <= 18'h20c00;\
    linear1_weight_array[6][68] <= 18'h00300;\
    linear1_weight_array[6][69] <= 18'h20080;\
    linear1_weight_array[6][70] <= 18'h00400;\
    linear1_weight_array[6][71] <= 18'h00600;\
    linear1_weight_array[6][72] <= 18'h20c00;\
    linear1_weight_array[6][73] <= 18'h00300;\
    linear1_weight_array[6][74] <= 18'h20080;\
    linear1_weight_array[6][75] <= 18'h00400;\
    linear1_weight_array[6][76] <= 18'h00600;\
    linear1_weight_array[6][77] <= 18'h20c00;\
    linear1_weight_array[6][78] <= 18'h00300;\
    linear1_weight_array[6][79] <= 18'h20080;\
    linear1_weight_array[6][80] <= 18'h00400;\
    linear1_weight_array[6][81] <= 18'h00600;\
    linear1_weight_array[6][82] <= 18'h20c00;\
    linear1_weight_array[6][83] <= 18'h00300;\
    linear1_weight_array[6][84] <= 18'h20080;\
    linear1_weight_array[6][85] <= 18'h00400;\
    linear1_weight_array[6][86] <= 18'h00600;\
    linear1_weight_array[6][87] <= 18'h20c00;\
    linear1_weight_array[6][88] <= 18'h00300;\
    linear1_weight_array[6][89] <= 18'h20080;\
    linear1_weight_array[6][90] <= 18'h00400;\
    linear1_weight_array[6][91] <= 18'h00600;\
    linear1_weight_array[6][92] <= 18'h20c00;\
    linear1_weight_array[6][93] <= 18'h00300;\
    linear1_weight_array[6][94] <= 18'h20080;\
    linear1_weight_array[6][95] <= 18'h00400;\
    linear1_weight_array[6][96] <= 18'h00600;\
    linear1_weight_array[6][97] <= 18'h20c00;\
    linear1_weight_array[6][98] <= 18'h00300;\
    linear1_weight_array[6][99] <= 18'h20080;\
    linear1_weight_array[6][100] <= 18'h00400;\
    linear1_weight_array[6][101] <= 18'h00600;\
    linear1_weight_array[6][102] <= 18'h20c00;\
    linear1_weight_array[6][103] <= 18'h00300;\
    linear1_weight_array[6][104] <= 18'h20080;\
    linear1_weight_array[6][105] <= 18'h00400;\
    linear1_weight_array[6][106] <= 18'h00600;\
    linear1_weight_array[6][107] <= 18'h20c00;\
    linear1_weight_array[6][108] <= 18'h00300;\
    linear1_weight_array[6][109] <= 18'h20080;\
    linear1_weight_array[6][110] <= 18'h00400;\
    linear1_weight_array[6][111] <= 18'h00600;\
    linear1_weight_array[6][112] <= 18'h20c00;\
    linear1_weight_array[6][113] <= 18'h00300;\
    linear1_weight_array[6][114] <= 18'h20080;\
    linear1_weight_array[6][115] <= 18'h00400;\
    linear1_weight_array[6][116] <= 18'h00600;\
    linear1_weight_array[6][117] <= 18'h20c00;\
    linear1_weight_array[6][118] <= 18'h00300;\
    linear1_weight_array[6][119] <= 18'h20080;\
    linear1_weight_array[6][120] <= 18'h00400;\
    linear1_weight_array[6][121] <= 18'h00600;\
    linear1_weight_array[6][122] <= 18'h20c00;\
    linear1_weight_array[6][123] <= 18'h00300;\
    linear1_weight_array[6][124] <= 18'h20080;\
    linear1_weight_array[6][125] <= 18'h00400;\
    linear1_weight_array[6][126] <= 18'h00600;\
    linear1_weight_array[6][127] <= 18'h20c00;\
    linear1_weight_array[6][128] <= 18'h00300;\
    linear1_weight_array[6][129] <= 18'h20080;\
    linear1_weight_array[6][130] <= 18'h00400;\
    linear1_weight_array[6][131] <= 18'h00600;\
    linear1_weight_array[6][132] <= 18'h20c00;\
    linear1_weight_array[6][133] <= 18'h00300;\
    linear1_weight_array[6][134] <= 18'h20080;\
    linear1_weight_array[6][135] <= 18'h00400;\
    linear1_weight_array[6][136] <= 18'h00600;\
    linear1_weight_array[6][137] <= 18'h20c00;\
    linear1_weight_array[6][138] <= 18'h00300;\
    linear1_weight_array[6][139] <= 18'h20080;\
    linear1_weight_array[6][140] <= 18'h00400;\
    linear1_weight_array[6][141] <= 18'h00600;\
    linear1_weight_array[6][142] <= 18'h20c00;\
    linear1_weight_array[6][143] <= 18'h00300;\
    linear1_weight_array[6][144] <= 18'h20080;\
    linear1_weight_array[6][145] <= 18'h00400;\
    linear1_weight_array[6][146] <= 18'h00600;\
    linear1_weight_array[6][147] <= 18'h20c00;\
    linear1_weight_array[6][148] <= 18'h00300;\
    linear1_weight_array[6][149] <= 18'h20080;\
    linear1_weight_array[7][0] <= 18'h00400;\
    linear1_weight_array[7][1] <= 18'h00600;\
    linear1_weight_array[7][2] <= 18'h20c00;\
    linear1_weight_array[7][3] <= 18'h00100;\
    linear1_weight_array[7][4] <= 18'h20080;\
    linear1_weight_array[7][5] <= 18'h00400;\
    linear1_weight_array[7][6] <= 18'h00600;\
    linear1_weight_array[7][7] <= 18'h20c00;\
    linear1_weight_array[7][8] <= 18'h00100;\
    linear1_weight_array[7][9] <= 18'h20080;\
    linear1_weight_array[7][10] <= 18'h00400;\
    linear1_weight_array[7][11] <= 18'h00600;\
    linear1_weight_array[7][12] <= 18'h20c00;\
    linear1_weight_array[7][13] <= 18'h00100;\
    linear1_weight_array[7][14] <= 18'h20080;\
    linear1_weight_array[7][15] <= 18'h00400;\
    linear1_weight_array[7][16] <= 18'h00600;\
    linear1_weight_array[7][17] <= 18'h20c00;\
    linear1_weight_array[7][18] <= 18'h00100;\
    linear1_weight_array[7][19] <= 18'h20080;\
    linear1_weight_array[7][20] <= 18'h00400;\
    linear1_weight_array[7][21] <= 18'h00600;\
    linear1_weight_array[7][22] <= 18'h20c00;\
    linear1_weight_array[7][23] <= 18'h00100;\
    linear1_weight_array[7][24] <= 18'h20080;\
    linear1_weight_array[7][25] <= 18'h00400;\
    linear1_weight_array[7][26] <= 18'h00600;\
    linear1_weight_array[7][27] <= 18'h20c00;\
    linear1_weight_array[7][28] <= 18'h00100;\
    linear1_weight_array[7][29] <= 18'h20080;\
    linear1_weight_array[7][30] <= 18'h00400;\
    linear1_weight_array[7][31] <= 18'h00600;\
    linear1_weight_array[7][32] <= 18'h20c00;\
    linear1_weight_array[7][33] <= 18'h00100;\
    linear1_weight_array[7][34] <= 18'h20080;\
    linear1_weight_array[7][35] <= 18'h00400;\
    linear1_weight_array[7][36] <= 18'h00600;\
    linear1_weight_array[7][37] <= 18'h20c00;\
    linear1_weight_array[7][38] <= 18'h00100;\
    linear1_weight_array[7][39] <= 18'h20080;\
    linear1_weight_array[7][40] <= 18'h00400;\
    linear1_weight_array[7][41] <= 18'h00600;\
    linear1_weight_array[7][42] <= 18'h20c00;\
    linear1_weight_array[7][43] <= 18'h00100;\
    linear1_weight_array[7][44] <= 18'h20080;\
    linear1_weight_array[7][45] <= 18'h00400;\
    linear1_weight_array[7][46] <= 18'h00600;\
    linear1_weight_array[7][47] <= 18'h20c00;\
    linear1_weight_array[7][48] <= 18'h00100;\
    linear1_weight_array[7][49] <= 18'h20080;\
    linear1_weight_array[7][50] <= 18'h00400;\
    linear1_weight_array[7][51] <= 18'h00600;\
    linear1_weight_array[7][52] <= 18'h20c00;\
    linear1_weight_array[7][53] <= 18'h00100;\
    linear1_weight_array[7][54] <= 18'h20080;\
    linear1_weight_array[7][55] <= 18'h00400;\
    linear1_weight_array[7][56] <= 18'h00600;\
    linear1_weight_array[7][57] <= 18'h20c00;\
    linear1_weight_array[7][58] <= 18'h00100;\
    linear1_weight_array[7][59] <= 18'h20080;\
    linear1_weight_array[7][60] <= 18'h00400;\
    linear1_weight_array[7][61] <= 18'h00600;\
    linear1_weight_array[7][62] <= 18'h20c00;\
    linear1_weight_array[7][63] <= 18'h00100;\
    linear1_weight_array[7][64] <= 18'h20080;\
    linear1_weight_array[7][65] <= 18'h00400;\
    linear1_weight_array[7][66] <= 18'h00600;\
    linear1_weight_array[7][67] <= 18'h20c00;\
    linear1_weight_array[7][68] <= 18'h00100;\
    linear1_weight_array[7][69] <= 18'h20080;\
    linear1_weight_array[7][70] <= 18'h00400;\
    linear1_weight_array[7][71] <= 18'h00600;\
    linear1_weight_array[7][72] <= 18'h20c00;\
    linear1_weight_array[7][73] <= 18'h00100;\
    linear1_weight_array[7][74] <= 18'h20080;\
    linear1_weight_array[7][75] <= 18'h00400;\
    linear1_weight_array[7][76] <= 18'h00600;\
    linear1_weight_array[7][77] <= 18'h20c00;\
    linear1_weight_array[7][78] <= 18'h00100;\
    linear1_weight_array[7][79] <= 18'h20080;\
    linear1_weight_array[7][80] <= 18'h00400;\
    linear1_weight_array[7][81] <= 18'h00600;\
    linear1_weight_array[7][82] <= 18'h20c00;\
    linear1_weight_array[7][83] <= 18'h00100;\
    linear1_weight_array[7][84] <= 18'h20080;\
    linear1_weight_array[7][85] <= 18'h00400;\
    linear1_weight_array[7][86] <= 18'h00600;\
    linear1_weight_array[7][87] <= 18'h20c00;\
    linear1_weight_array[7][88] <= 18'h00100;\
    linear1_weight_array[7][89] <= 18'h20080;\
    linear1_weight_array[7][90] <= 18'h00400;\
    linear1_weight_array[7][91] <= 18'h00600;\
    linear1_weight_array[7][92] <= 18'h20c00;\
    linear1_weight_array[7][93] <= 18'h00100;\
    linear1_weight_array[7][94] <= 18'h20080;\
    linear1_weight_array[7][95] <= 18'h00400;\
    linear1_weight_array[7][96] <= 18'h00600;\
    linear1_weight_array[7][97] <= 18'h20c00;\
    linear1_weight_array[7][98] <= 18'h00100;\
    linear1_weight_array[7][99] <= 18'h20080;\
    linear1_weight_array[7][100] <= 18'h00400;\
    linear1_weight_array[7][101] <= 18'h00600;\
    linear1_weight_array[7][102] <= 18'h20c00;\
    linear1_weight_array[7][103] <= 18'h00100;\
    linear1_weight_array[7][104] <= 18'h20080;\
    linear1_weight_array[7][105] <= 18'h00400;\
    linear1_weight_array[7][106] <= 18'h00600;\
    linear1_weight_array[7][107] <= 18'h20c00;\
    linear1_weight_array[7][108] <= 18'h00100;\
    linear1_weight_array[7][109] <= 18'h20080;\
    linear1_weight_array[7][110] <= 18'h00400;\
    linear1_weight_array[7][111] <= 18'h00600;\
    linear1_weight_array[7][112] <= 18'h20c00;\
    linear1_weight_array[7][113] <= 18'h00100;\
    linear1_weight_array[7][114] <= 18'h20080;\
    linear1_weight_array[7][115] <= 18'h00400;\
    linear1_weight_array[7][116] <= 18'h00600;\
    linear1_weight_array[7][117] <= 18'h20c00;\
    linear1_weight_array[7][118] <= 18'h00100;\
    linear1_weight_array[7][119] <= 18'h20080;\
    linear1_weight_array[7][120] <= 18'h00400;\
    linear1_weight_array[7][121] <= 18'h00600;\
    linear1_weight_array[7][122] <= 18'h20c00;\
    linear1_weight_array[7][123] <= 18'h00100;\
    linear1_weight_array[7][124] <= 18'h20080;\
    linear1_weight_array[7][125] <= 18'h00400;\
    linear1_weight_array[7][126] <= 18'h00600;\
    linear1_weight_array[7][127] <= 18'h20c00;\
    linear1_weight_array[7][128] <= 18'h00100;\
    linear1_weight_array[7][129] <= 18'h20080;\
    linear1_weight_array[7][130] <= 18'h00400;\
    linear1_weight_array[7][131] <= 18'h00600;\
    linear1_weight_array[7][132] <= 18'h20c00;\
    linear1_weight_array[7][133] <= 18'h00100;\
    linear1_weight_array[7][134] <= 18'h20080;\
    linear1_weight_array[7][135] <= 18'h00400;\
    linear1_weight_array[7][136] <= 18'h00600;\
    linear1_weight_array[7][137] <= 18'h20c00;\
    linear1_weight_array[7][138] <= 18'h00100;\
    linear1_weight_array[7][139] <= 18'h20080;\
    linear1_weight_array[7][140] <= 18'h00400;\
    linear1_weight_array[7][141] <= 18'h00600;\
    linear1_weight_array[7][142] <= 18'h20c00;\
    linear1_weight_array[7][143] <= 18'h00100;\
    linear1_weight_array[7][144] <= 18'h20080;\
    linear1_weight_array[7][145] <= 18'h00400;\
    linear1_weight_array[7][146] <= 18'h00600;\
    linear1_weight_array[7][147] <= 18'h20c00;\
    linear1_weight_array[7][148] <= 18'h00100;\
    linear1_weight_array[7][149] <= 18'h20080;\
    linear1_weight_array[8][0] <= 18'h00400;\
    linear1_weight_array[8][1] <= 18'h00600;\
    linear1_weight_array[8][2] <= 18'h20c00;\
    linear1_weight_array[8][3] <= 18'h00300;\
    linear1_weight_array[8][4] <= 18'h20080;\
    linear1_weight_array[8][5] <= 18'h00400;\
    linear1_weight_array[8][6] <= 18'h00600;\
    linear1_weight_array[8][7] <= 18'h20c00;\
    linear1_weight_array[8][8] <= 18'h00300;\
    linear1_weight_array[8][9] <= 18'h20080;\
    linear1_weight_array[8][10] <= 18'h00400;\
    linear1_weight_array[8][11] <= 18'h00600;\
    linear1_weight_array[8][12] <= 18'h20c00;\
    linear1_weight_array[8][13] <= 18'h00300;\
    linear1_weight_array[8][14] <= 18'h20080;\
    linear1_weight_array[8][15] <= 18'h00400;\
    linear1_weight_array[8][16] <= 18'h00600;\
    linear1_weight_array[8][17] <= 18'h20c00;\
    linear1_weight_array[8][18] <= 18'h00300;\
    linear1_weight_array[8][19] <= 18'h20080;\
    linear1_weight_array[8][20] <= 18'h00400;\
    linear1_weight_array[8][21] <= 18'h00600;\
    linear1_weight_array[8][22] <= 18'h20c00;\
    linear1_weight_array[8][23] <= 18'h00300;\
    linear1_weight_array[8][24] <= 18'h20080;\
    linear1_weight_array[8][25] <= 18'h00400;\
    linear1_weight_array[8][26] <= 18'h00600;\
    linear1_weight_array[8][27] <= 18'h20c00;\
    linear1_weight_array[8][28] <= 18'h00300;\
    linear1_weight_array[8][29] <= 18'h20080;\
    linear1_weight_array[8][30] <= 18'h00400;\
    linear1_weight_array[8][31] <= 18'h00600;\
    linear1_weight_array[8][32] <= 18'h20c00;\
    linear1_weight_array[8][33] <= 18'h00300;\
    linear1_weight_array[8][34] <= 18'h20080;\
    linear1_weight_array[8][35] <= 18'h00400;\
    linear1_weight_array[8][36] <= 18'h00600;\
    linear1_weight_array[8][37] <= 18'h20c00;\
    linear1_weight_array[8][38] <= 18'h00300;\
    linear1_weight_array[8][39] <= 18'h20080;\
    linear1_weight_array[8][40] <= 18'h00400;\
    linear1_weight_array[8][41] <= 18'h00600;\
    linear1_weight_array[8][42] <= 18'h20c00;\
    linear1_weight_array[8][43] <= 18'h00300;\
    linear1_weight_array[8][44] <= 18'h20080;\
    linear1_weight_array[8][45] <= 18'h00400;\
    linear1_weight_array[8][46] <= 18'h00600;\
    linear1_weight_array[8][47] <= 18'h20c00;\
    linear1_weight_array[8][48] <= 18'h00300;\
    linear1_weight_array[8][49] <= 18'h20080;\
    linear1_weight_array[8][50] <= 18'h00400;\
    linear1_weight_array[8][51] <= 18'h00600;\
    linear1_weight_array[8][52] <= 18'h20c00;\
    linear1_weight_array[8][53] <= 18'h00300;\
    linear1_weight_array[8][54] <= 18'h20080;\
    linear1_weight_array[8][55] <= 18'h00400;\
    linear1_weight_array[8][56] <= 18'h00600;\
    linear1_weight_array[8][57] <= 18'h20c00;\
    linear1_weight_array[8][58] <= 18'h00300;\
    linear1_weight_array[8][59] <= 18'h20080;\
    linear1_weight_array[8][60] <= 18'h00400;\
    linear1_weight_array[8][61] <= 18'h00600;\
    linear1_weight_array[8][62] <= 18'h20c00;\
    linear1_weight_array[8][63] <= 18'h00300;\
    linear1_weight_array[8][64] <= 18'h20080;\
    linear1_weight_array[8][65] <= 18'h00400;\
    linear1_weight_array[8][66] <= 18'h00600;\
    linear1_weight_array[8][67] <= 18'h20c00;\
    linear1_weight_array[8][68] <= 18'h00300;\
    linear1_weight_array[8][69] <= 18'h20080;\
    linear1_weight_array[8][70] <= 18'h00400;\
    linear1_weight_array[8][71] <= 18'h00600;\
    linear1_weight_array[8][72] <= 18'h20c00;\
    linear1_weight_array[8][73] <= 18'h00300;\
    linear1_weight_array[8][74] <= 18'h20080;\
    linear1_weight_array[8][75] <= 18'h00400;\
    linear1_weight_array[8][76] <= 18'h00600;\
    linear1_weight_array[8][77] <= 18'h20c00;\
    linear1_weight_array[8][78] <= 18'h00300;\
    linear1_weight_array[8][79] <= 18'h20080;\
    linear1_weight_array[8][80] <= 18'h00400;\
    linear1_weight_array[8][81] <= 18'h00600;\
    linear1_weight_array[8][82] <= 18'h20c00;\
    linear1_weight_array[8][83] <= 18'h00300;\
    linear1_weight_array[8][84] <= 18'h20080;\
    linear1_weight_array[8][85] <= 18'h00400;\
    linear1_weight_array[8][86] <= 18'h00600;\
    linear1_weight_array[8][87] <= 18'h20c00;\
    linear1_weight_array[8][88] <= 18'h00300;\
    linear1_weight_array[8][89] <= 18'h20080;\
    linear1_weight_array[8][90] <= 18'h00400;\
    linear1_weight_array[8][91] <= 18'h00600;\
    linear1_weight_array[8][92] <= 18'h20c00;\
    linear1_weight_array[8][93] <= 18'h00300;\
    linear1_weight_array[8][94] <= 18'h20080;\
    linear1_weight_array[8][95] <= 18'h00400;\
    linear1_weight_array[8][96] <= 18'h00600;\
    linear1_weight_array[8][97] <= 18'h20c00;\
    linear1_weight_array[8][98] <= 18'h00300;\
    linear1_weight_array[8][99] <= 18'h20080;\
    linear1_weight_array[8][100] <= 18'h00400;\
    linear1_weight_array[8][101] <= 18'h00600;\
    linear1_weight_array[8][102] <= 18'h20c00;\
    linear1_weight_array[8][103] <= 18'h00300;\
    linear1_weight_array[8][104] <= 18'h20080;\
    linear1_weight_array[8][105] <= 18'h00400;\
    linear1_weight_array[8][106] <= 18'h00600;\
    linear1_weight_array[8][107] <= 18'h20c00;\
    linear1_weight_array[8][108] <= 18'h00300;\
    linear1_weight_array[8][109] <= 18'h20080;\
    linear1_weight_array[8][110] <= 18'h00400;\
    linear1_weight_array[8][111] <= 18'h00600;\
    linear1_weight_array[8][112] <= 18'h20c00;\
    linear1_weight_array[8][113] <= 18'h00300;\
    linear1_weight_array[8][114] <= 18'h20080;\
    linear1_weight_array[8][115] <= 18'h00400;\
    linear1_weight_array[8][116] <= 18'h00600;\
    linear1_weight_array[8][117] <= 18'h20c00;\
    linear1_weight_array[8][118] <= 18'h00300;\
    linear1_weight_array[8][119] <= 18'h20080;\
    linear1_weight_array[8][120] <= 18'h00400;\
    linear1_weight_array[8][121] <= 18'h00600;\
    linear1_weight_array[8][122] <= 18'h20c00;\
    linear1_weight_array[8][123] <= 18'h00300;\
    linear1_weight_array[8][124] <= 18'h20080;\
    linear1_weight_array[8][125] <= 18'h00400;\
    linear1_weight_array[8][126] <= 18'h00600;\
    linear1_weight_array[8][127] <= 18'h20c00;\
    linear1_weight_array[8][128] <= 18'h00300;\
    linear1_weight_array[8][129] <= 18'h20080;\
    linear1_weight_array[8][130] <= 18'h00400;\
    linear1_weight_array[8][131] <= 18'h00600;\
    linear1_weight_array[8][132] <= 18'h20c00;\
    linear1_weight_array[8][133] <= 18'h00300;\
    linear1_weight_array[8][134] <= 18'h20080;\
    linear1_weight_array[8][135] <= 18'h00400;\
    linear1_weight_array[8][136] <= 18'h00600;\
    linear1_weight_array[8][137] <= 18'h20c00;\
    linear1_weight_array[8][138] <= 18'h00300;\
    linear1_weight_array[8][139] <= 18'h20080;\
    linear1_weight_array[8][140] <= 18'h00400;\
    linear1_weight_array[8][141] <= 18'h00600;\
    linear1_weight_array[8][142] <= 18'h20c00;\
    linear1_weight_array[8][143] <= 18'h00300;\
    linear1_weight_array[8][144] <= 18'h20080;\
    linear1_weight_array[8][145] <= 18'h00400;\
    linear1_weight_array[8][146] <= 18'h00600;\
    linear1_weight_array[8][147] <= 18'h20c00;\
    linear1_weight_array[8][148] <= 18'h00300;\
    linear1_weight_array[8][149] <= 18'h20080;\
    linear1_weight_array[9][0] <= 18'h00400;\
    linear1_weight_array[9][1] <= 18'h00600;\
    linear1_weight_array[9][2] <= 18'h20c00;\
    linear1_weight_array[9][3] <= 18'h00100;\
    linear1_weight_array[9][4] <= 18'h20080;\
    linear1_weight_array[9][5] <= 18'h00400;\
    linear1_weight_array[9][6] <= 18'h00600;\
    linear1_weight_array[9][7] <= 18'h20c00;\
    linear1_weight_array[9][8] <= 18'h00100;\
    linear1_weight_array[9][9] <= 18'h20080;\
    linear1_weight_array[9][10] <= 18'h00400;\
    linear1_weight_array[9][11] <= 18'h00600;\
    linear1_weight_array[9][12] <= 18'h20c00;\
    linear1_weight_array[9][13] <= 18'h00100;\
    linear1_weight_array[9][14] <= 18'h20080;\
    linear1_weight_array[9][15] <= 18'h00400;\
    linear1_weight_array[9][16] <= 18'h00600;\
    linear1_weight_array[9][17] <= 18'h20c00;\
    linear1_weight_array[9][18] <= 18'h00100;\
    linear1_weight_array[9][19] <= 18'h20080;\
    linear1_weight_array[9][20] <= 18'h00400;\
    linear1_weight_array[9][21] <= 18'h00600;\
    linear1_weight_array[9][22] <= 18'h20c00;\
    linear1_weight_array[9][23] <= 18'h00100;\
    linear1_weight_array[9][24] <= 18'h20080;\
    linear1_weight_array[9][25] <= 18'h00400;\
    linear1_weight_array[9][26] <= 18'h00600;\
    linear1_weight_array[9][27] <= 18'h20c00;\
    linear1_weight_array[9][28] <= 18'h00100;\
    linear1_weight_array[9][29] <= 18'h20080;\
    linear1_weight_array[9][30] <= 18'h00400;\
    linear1_weight_array[9][31] <= 18'h00600;\
    linear1_weight_array[9][32] <= 18'h20c00;\
    linear1_weight_array[9][33] <= 18'h00100;\
    linear1_weight_array[9][34] <= 18'h20080;\
    linear1_weight_array[9][35] <= 18'h00400;\
    linear1_weight_array[9][36] <= 18'h00600;\
    linear1_weight_array[9][37] <= 18'h20c00;\
    linear1_weight_array[9][38] <= 18'h00100;\
    linear1_weight_array[9][39] <= 18'h20080;\
    linear1_weight_array[9][40] <= 18'h00400;\
    linear1_weight_array[9][41] <= 18'h00600;\
    linear1_weight_array[9][42] <= 18'h20c00;\
    linear1_weight_array[9][43] <= 18'h00100;\
    linear1_weight_array[9][44] <= 18'h20080;\
    linear1_weight_array[9][45] <= 18'h00400;\
    linear1_weight_array[9][46] <= 18'h00600;\
    linear1_weight_array[9][47] <= 18'h20c00;\
    linear1_weight_array[9][48] <= 18'h00100;\
    linear1_weight_array[9][49] <= 18'h20080;\
    linear1_weight_array[9][50] <= 18'h00400;\
    linear1_weight_array[9][51] <= 18'h00600;\
    linear1_weight_array[9][52] <= 18'h20c00;\
    linear1_weight_array[9][53] <= 18'h00100;\
    linear1_weight_array[9][54] <= 18'h20080;\
    linear1_weight_array[9][55] <= 18'h00400;\
    linear1_weight_array[9][56] <= 18'h00600;\
    linear1_weight_array[9][57] <= 18'h20c00;\
    linear1_weight_array[9][58] <= 18'h00100;\
    linear1_weight_array[9][59] <= 18'h20080;\
    linear1_weight_array[9][60] <= 18'h00400;\
    linear1_weight_array[9][61] <= 18'h00600;\
    linear1_weight_array[9][62] <= 18'h20c00;\
    linear1_weight_array[9][63] <= 18'h00100;\
    linear1_weight_array[9][64] <= 18'h20080;\
    linear1_weight_array[9][65] <= 18'h00400;\
    linear1_weight_array[9][66] <= 18'h00600;\
    linear1_weight_array[9][67] <= 18'h20c00;\
    linear1_weight_array[9][68] <= 18'h00100;\
    linear1_weight_array[9][69] <= 18'h20080;\
    linear1_weight_array[9][70] <= 18'h00400;\
    linear1_weight_array[9][71] <= 18'h00600;\
    linear1_weight_array[9][72] <= 18'h20c00;\
    linear1_weight_array[9][73] <= 18'h00100;\
    linear1_weight_array[9][74] <= 18'h20080;\
    linear1_weight_array[9][75] <= 18'h00400;\
    linear1_weight_array[9][76] <= 18'h00600;\
    linear1_weight_array[9][77] <= 18'h20c00;\
    linear1_weight_array[9][78] <= 18'h00100;\
    linear1_weight_array[9][79] <= 18'h20080;\
    linear1_weight_array[9][80] <= 18'h00400;\
    linear1_weight_array[9][81] <= 18'h00600;\
    linear1_weight_array[9][82] <= 18'h20c00;\
    linear1_weight_array[9][83] <= 18'h00100;\
    linear1_weight_array[9][84] <= 18'h20080;\
    linear1_weight_array[9][85] <= 18'h00400;\
    linear1_weight_array[9][86] <= 18'h00600;\
    linear1_weight_array[9][87] <= 18'h20c00;\
    linear1_weight_array[9][88] <= 18'h00100;\
    linear1_weight_array[9][89] <= 18'h20080;\
    linear1_weight_array[9][90] <= 18'h00400;\
    linear1_weight_array[9][91] <= 18'h00600;\
    linear1_weight_array[9][92] <= 18'h20c00;\
    linear1_weight_array[9][93] <= 18'h00100;\
    linear1_weight_array[9][94] <= 18'h20080;\
    linear1_weight_array[9][95] <= 18'h00400;\
    linear1_weight_array[9][96] <= 18'h00600;\
    linear1_weight_array[9][97] <= 18'h20c00;\
    linear1_weight_array[9][98] <= 18'h00100;\
    linear1_weight_array[9][99] <= 18'h20080;\
    linear1_weight_array[9][100] <= 18'h00400;\
    linear1_weight_array[9][101] <= 18'h00600;\
    linear1_weight_array[9][102] <= 18'h20c00;\
    linear1_weight_array[9][103] <= 18'h00100;\
    linear1_weight_array[9][104] <= 18'h20080;\
    linear1_weight_array[9][105] <= 18'h00400;\
    linear1_weight_array[9][106] <= 18'h00600;\
    linear1_weight_array[9][107] <= 18'h20c00;\
    linear1_weight_array[9][108] <= 18'h00100;\
    linear1_weight_array[9][109] <= 18'h20080;\
    linear1_weight_array[9][110] <= 18'h00400;\
    linear1_weight_array[9][111] <= 18'h00600;\
    linear1_weight_array[9][112] <= 18'h20c00;\
    linear1_weight_array[9][113] <= 18'h00100;\
    linear1_weight_array[9][114] <= 18'h20080;\
    linear1_weight_array[9][115] <= 18'h00400;\
    linear1_weight_array[9][116] <= 18'h00600;\
    linear1_weight_array[9][117] <= 18'h20c00;\
    linear1_weight_array[9][118] <= 18'h00100;\
    linear1_weight_array[9][119] <= 18'h20080;\
    linear1_weight_array[9][120] <= 18'h00400;\
    linear1_weight_array[9][121] <= 18'h00600;\
    linear1_weight_array[9][122] <= 18'h20c00;\
    linear1_weight_array[9][123] <= 18'h00100;\
    linear1_weight_array[9][124] <= 18'h20080;\
    linear1_weight_array[9][125] <= 18'h00400;\
    linear1_weight_array[9][126] <= 18'h00600;\
    linear1_weight_array[9][127] <= 18'h20c00;\
    linear1_weight_array[9][128] <= 18'h00100;\
    linear1_weight_array[9][129] <= 18'h20080;\
    linear1_weight_array[9][130] <= 18'h00400;\
    linear1_weight_array[9][131] <= 18'h00600;\
    linear1_weight_array[9][132] <= 18'h20c00;\
    linear1_weight_array[9][133] <= 18'h00100;\
    linear1_weight_array[9][134] <= 18'h20080;\
    linear1_weight_array[9][135] <= 18'h00400;\
    linear1_weight_array[9][136] <= 18'h00600;\
    linear1_weight_array[9][137] <= 18'h20c00;\
    linear1_weight_array[9][138] <= 18'h00100;\
    linear1_weight_array[9][139] <= 18'h20080;\
    linear1_weight_array[9][140] <= 18'h00400;\
    linear1_weight_array[9][141] <= 18'h00600;\
    linear1_weight_array[9][142] <= 18'h20c00;\
    linear1_weight_array[9][143] <= 18'h00100;\
    linear1_weight_array[9][144] <= 18'h20080;\
    linear1_weight_array[9][145] <= 18'h00400;\
    linear1_weight_array[9][146] <= 18'h00600;\
    linear1_weight_array[9][147] <= 18'h20c00;\
    linear1_weight_array[9][148] <= 18'h00100;\
    linear1_weight_array[9][149] <= 18'h20080;\
    linear1_weight_array[10][0] <= 18'h00400;\
    linear1_weight_array[10][1] <= 18'h00600;\
    linear1_weight_array[10][2] <= 18'h20c00;\
    linear1_weight_array[10][3] <= 18'h00300;\
    linear1_weight_array[10][4] <= 18'h20080;\
    linear1_weight_array[10][5] <= 18'h00400;\
    linear1_weight_array[10][6] <= 18'h00600;\
    linear1_weight_array[10][7] <= 18'h20c00;\
    linear1_weight_array[10][8] <= 18'h00300;\
    linear1_weight_array[10][9] <= 18'h20080;\
    linear1_weight_array[10][10] <= 18'h00400;\
    linear1_weight_array[10][11] <= 18'h00600;\
    linear1_weight_array[10][12] <= 18'h20c00;\
    linear1_weight_array[10][13] <= 18'h00300;\
    linear1_weight_array[10][14] <= 18'h20080;\
    linear1_weight_array[10][15] <= 18'h00400;\
    linear1_weight_array[10][16] <= 18'h00600;\
    linear1_weight_array[10][17] <= 18'h20c00;\
    linear1_weight_array[10][18] <= 18'h00300;\
    linear1_weight_array[10][19] <= 18'h20080;\
    linear1_weight_array[10][20] <= 18'h00400;\
    linear1_weight_array[10][21] <= 18'h00600;\
    linear1_weight_array[10][22] <= 18'h20c00;\
    linear1_weight_array[10][23] <= 18'h00300;\
    linear1_weight_array[10][24] <= 18'h20080;\
    linear1_weight_array[10][25] <= 18'h00400;\
    linear1_weight_array[10][26] <= 18'h00600;\
    linear1_weight_array[10][27] <= 18'h20c00;\
    linear1_weight_array[10][28] <= 18'h00300;\
    linear1_weight_array[10][29] <= 18'h20080;\
    linear1_weight_array[10][30] <= 18'h00400;\
    linear1_weight_array[10][31] <= 18'h00600;\
    linear1_weight_array[10][32] <= 18'h20c00;\
    linear1_weight_array[10][33] <= 18'h00300;\
    linear1_weight_array[10][34] <= 18'h20080;\
    linear1_weight_array[10][35] <= 18'h00400;\
    linear1_weight_array[10][36] <= 18'h00600;\
    linear1_weight_array[10][37] <= 18'h20c00;\
    linear1_weight_array[10][38] <= 18'h00300;\
    linear1_weight_array[10][39] <= 18'h20080;\
    linear1_weight_array[10][40] <= 18'h00400;\
    linear1_weight_array[10][41] <= 18'h00600;\
    linear1_weight_array[10][42] <= 18'h20c00;\
    linear1_weight_array[10][43] <= 18'h00300;\
    linear1_weight_array[10][44] <= 18'h20080;\
    linear1_weight_array[10][45] <= 18'h00400;\
    linear1_weight_array[10][46] <= 18'h00600;\
    linear1_weight_array[10][47] <= 18'h20c00;\
    linear1_weight_array[10][48] <= 18'h00300;\
    linear1_weight_array[10][49] <= 18'h20080;\
    linear1_weight_array[10][50] <= 18'h00400;\
    linear1_weight_array[10][51] <= 18'h00600;\
    linear1_weight_array[10][52] <= 18'h20c00;\
    linear1_weight_array[10][53] <= 18'h00300;\
    linear1_weight_array[10][54] <= 18'h20080;\
    linear1_weight_array[10][55] <= 18'h00400;\
    linear1_weight_array[10][56] <= 18'h00600;\
    linear1_weight_array[10][57] <= 18'h20c00;\
    linear1_weight_array[10][58] <= 18'h00300;\
    linear1_weight_array[10][59] <= 18'h20080;\
    linear1_weight_array[10][60] <= 18'h00400;\
    linear1_weight_array[10][61] <= 18'h00600;\
    linear1_weight_array[10][62] <= 18'h20c00;\
    linear1_weight_array[10][63] <= 18'h00300;\
    linear1_weight_array[10][64] <= 18'h20080;\
    linear1_weight_array[10][65] <= 18'h00400;\
    linear1_weight_array[10][66] <= 18'h00600;\
    linear1_weight_array[10][67] <= 18'h20c00;\
    linear1_weight_array[10][68] <= 18'h00300;\
    linear1_weight_array[10][69] <= 18'h20080;\
    linear1_weight_array[10][70] <= 18'h00400;\
    linear1_weight_array[10][71] <= 18'h00600;\
    linear1_weight_array[10][72] <= 18'h20c00;\
    linear1_weight_array[10][73] <= 18'h00300;\
    linear1_weight_array[10][74] <= 18'h20080;\
    linear1_weight_array[10][75] <= 18'h00400;\
    linear1_weight_array[10][76] <= 18'h00600;\
    linear1_weight_array[10][77] <= 18'h20c00;\
    linear1_weight_array[10][78] <= 18'h00300;\
    linear1_weight_array[10][79] <= 18'h20080;\
    linear1_weight_array[10][80] <= 18'h00400;\
    linear1_weight_array[10][81] <= 18'h00600;\
    linear1_weight_array[10][82] <= 18'h20c00;\
    linear1_weight_array[10][83] <= 18'h00300;\
    linear1_weight_array[10][84] <= 18'h20080;\
    linear1_weight_array[10][85] <= 18'h00400;\
    linear1_weight_array[10][86] <= 18'h00600;\
    linear1_weight_array[10][87] <= 18'h20c00;\
    linear1_weight_array[10][88] <= 18'h00300;\
    linear1_weight_array[10][89] <= 18'h20080;\
    linear1_weight_array[10][90] <= 18'h00400;\
    linear1_weight_array[10][91] <= 18'h00600;\
    linear1_weight_array[10][92] <= 18'h20c00;\
    linear1_weight_array[10][93] <= 18'h00300;\
    linear1_weight_array[10][94] <= 18'h20080;\
    linear1_weight_array[10][95] <= 18'h00400;\
    linear1_weight_array[10][96] <= 18'h00600;\
    linear1_weight_array[10][97] <= 18'h20c00;\
    linear1_weight_array[10][98] <= 18'h00300;\
    linear1_weight_array[10][99] <= 18'h20080;\
    linear1_weight_array[10][100] <= 18'h00400;\
    linear1_weight_array[10][101] <= 18'h00600;\
    linear1_weight_array[10][102] <= 18'h20c00;\
    linear1_weight_array[10][103] <= 18'h00300;\
    linear1_weight_array[10][104] <= 18'h20080;\
    linear1_weight_array[10][105] <= 18'h00400;\
    linear1_weight_array[10][106] <= 18'h00600;\
    linear1_weight_array[10][107] <= 18'h20c00;\
    linear1_weight_array[10][108] <= 18'h00300;\
    linear1_weight_array[10][109] <= 18'h20080;\
    linear1_weight_array[10][110] <= 18'h00400;\
    linear1_weight_array[10][111] <= 18'h00600;\
    linear1_weight_array[10][112] <= 18'h20c00;\
    linear1_weight_array[10][113] <= 18'h00300;\
    linear1_weight_array[10][114] <= 18'h20080;\
    linear1_weight_array[10][115] <= 18'h00400;\
    linear1_weight_array[10][116] <= 18'h00600;\
    linear1_weight_array[10][117] <= 18'h20c00;\
    linear1_weight_array[10][118] <= 18'h00300;\
    linear1_weight_array[10][119] <= 18'h20080;\
    linear1_weight_array[10][120] <= 18'h00400;\
    linear1_weight_array[10][121] <= 18'h00600;\
    linear1_weight_array[10][122] <= 18'h20c00;\
    linear1_weight_array[10][123] <= 18'h00300;\
    linear1_weight_array[10][124] <= 18'h20080;\
    linear1_weight_array[10][125] <= 18'h00400;\
    linear1_weight_array[10][126] <= 18'h00600;\
    linear1_weight_array[10][127] <= 18'h20c00;\
    linear1_weight_array[10][128] <= 18'h00300;\
    linear1_weight_array[10][129] <= 18'h20080;\
    linear1_weight_array[10][130] <= 18'h00400;\
    linear1_weight_array[10][131] <= 18'h00600;\
    linear1_weight_array[10][132] <= 18'h20c00;\
    linear1_weight_array[10][133] <= 18'h00300;\
    linear1_weight_array[10][134] <= 18'h20080;\
    linear1_weight_array[10][135] <= 18'h00400;\
    linear1_weight_array[10][136] <= 18'h00600;\
    linear1_weight_array[10][137] <= 18'h20c00;\
    linear1_weight_array[10][138] <= 18'h00300;\
    linear1_weight_array[10][139] <= 18'h20080;\
    linear1_weight_array[10][140] <= 18'h00400;\
    linear1_weight_array[10][141] <= 18'h00600;\
    linear1_weight_array[10][142] <= 18'h20c00;\
    linear1_weight_array[10][143] <= 18'h00300;\
    linear1_weight_array[10][144] <= 18'h20080;\
    linear1_weight_array[10][145] <= 18'h00400;\
    linear1_weight_array[10][146] <= 18'h00600;\
    linear1_weight_array[10][147] <= 18'h20c00;\
    linear1_weight_array[10][148] <= 18'h00300;\
    linear1_weight_array[10][149] <= 18'h20080;\
    linear1_weight_array[11][0] <= 18'h00400;\
    linear1_weight_array[11][1] <= 18'h00600;\
    linear1_weight_array[11][2] <= 18'h20c00;\
    linear1_weight_array[11][3] <= 18'h00100;\
    linear1_weight_array[11][4] <= 18'h20080;\
    linear1_weight_array[11][5] <= 18'h00400;\
    linear1_weight_array[11][6] <= 18'h00600;\
    linear1_weight_array[11][7] <= 18'h20c00;\
    linear1_weight_array[11][8] <= 18'h00100;\
    linear1_weight_array[11][9] <= 18'h20080;\
    linear1_weight_array[11][10] <= 18'h00400;\
    linear1_weight_array[11][11] <= 18'h00600;\
    linear1_weight_array[11][12] <= 18'h20c00;\
    linear1_weight_array[11][13] <= 18'h00100;\
    linear1_weight_array[11][14] <= 18'h20080;\
    linear1_weight_array[11][15] <= 18'h00400;\
    linear1_weight_array[11][16] <= 18'h00600;\
    linear1_weight_array[11][17] <= 18'h20c00;\
    linear1_weight_array[11][18] <= 18'h00100;\
    linear1_weight_array[11][19] <= 18'h20080;\
    linear1_weight_array[11][20] <= 18'h00400;\
    linear1_weight_array[11][21] <= 18'h00600;\
    linear1_weight_array[11][22] <= 18'h20c00;\
    linear1_weight_array[11][23] <= 18'h00100;\
    linear1_weight_array[11][24] <= 18'h20080;\
    linear1_weight_array[11][25] <= 18'h00400;\
    linear1_weight_array[11][26] <= 18'h00600;\
    linear1_weight_array[11][27] <= 18'h20c00;\
    linear1_weight_array[11][28] <= 18'h00100;\
    linear1_weight_array[11][29] <= 18'h20080;\
    linear1_weight_array[11][30] <= 18'h00400;\
    linear1_weight_array[11][31] <= 18'h00600;\
    linear1_weight_array[11][32] <= 18'h20c00;\
    linear1_weight_array[11][33] <= 18'h00100;\
    linear1_weight_array[11][34] <= 18'h20080;\
    linear1_weight_array[11][35] <= 18'h00400;\
    linear1_weight_array[11][36] <= 18'h00600;\
    linear1_weight_array[11][37] <= 18'h20c00;\
    linear1_weight_array[11][38] <= 18'h00100;\
    linear1_weight_array[11][39] <= 18'h20080;\
    linear1_weight_array[11][40] <= 18'h00400;\
    linear1_weight_array[11][41] <= 18'h00600;\
    linear1_weight_array[11][42] <= 18'h20c00;\
    linear1_weight_array[11][43] <= 18'h00100;\
    linear1_weight_array[11][44] <= 18'h20080;\
    linear1_weight_array[11][45] <= 18'h00400;\
    linear1_weight_array[11][46] <= 18'h00600;\
    linear1_weight_array[11][47] <= 18'h20c00;\
    linear1_weight_array[11][48] <= 18'h00100;\
    linear1_weight_array[11][49] <= 18'h20080;\
    linear1_weight_array[11][50] <= 18'h00400;\
    linear1_weight_array[11][51] <= 18'h00600;\
    linear1_weight_array[11][52] <= 18'h20c00;\
    linear1_weight_array[11][53] <= 18'h00100;\
    linear1_weight_array[11][54] <= 18'h20080;\
    linear1_weight_array[11][55] <= 18'h00400;\
    linear1_weight_array[11][56] <= 18'h00600;\
    linear1_weight_array[11][57] <= 18'h20c00;\
    linear1_weight_array[11][58] <= 18'h00100;\
    linear1_weight_array[11][59] <= 18'h20080;\
    linear1_weight_array[11][60] <= 18'h00400;\
    linear1_weight_array[11][61] <= 18'h00600;\
    linear1_weight_array[11][62] <= 18'h20c00;\
    linear1_weight_array[11][63] <= 18'h00100;\
    linear1_weight_array[11][64] <= 18'h20080;\
    linear1_weight_array[11][65] <= 18'h00400;\
    linear1_weight_array[11][66] <= 18'h00600;\
    linear1_weight_array[11][67] <= 18'h20c00;\
    linear1_weight_array[11][68] <= 18'h00100;\
    linear1_weight_array[11][69] <= 18'h20080;\
    linear1_weight_array[11][70] <= 18'h00400;\
    linear1_weight_array[11][71] <= 18'h00600;\
    linear1_weight_array[11][72] <= 18'h20c00;\
    linear1_weight_array[11][73] <= 18'h00100;\
    linear1_weight_array[11][74] <= 18'h20080;\
    linear1_weight_array[11][75] <= 18'h00400;\
    linear1_weight_array[11][76] <= 18'h00600;\
    linear1_weight_array[11][77] <= 18'h20c00;\
    linear1_weight_array[11][78] <= 18'h00100;\
    linear1_weight_array[11][79] <= 18'h20080;\
    linear1_weight_array[11][80] <= 18'h00400;\
    linear1_weight_array[11][81] <= 18'h00600;\
    linear1_weight_array[11][82] <= 18'h20c00;\
    linear1_weight_array[11][83] <= 18'h00100;\
    linear1_weight_array[11][84] <= 18'h20080;\
    linear1_weight_array[11][85] <= 18'h00400;\
    linear1_weight_array[11][86] <= 18'h00600;\
    linear1_weight_array[11][87] <= 18'h20c00;\
    linear1_weight_array[11][88] <= 18'h00100;\
    linear1_weight_array[11][89] <= 18'h20080;\
    linear1_weight_array[11][90] <= 18'h00400;\
    linear1_weight_array[11][91] <= 18'h00600;\
    linear1_weight_array[11][92] <= 18'h20c00;\
    linear1_weight_array[11][93] <= 18'h00100;\
    linear1_weight_array[11][94] <= 18'h20080;\
    linear1_weight_array[11][95] <= 18'h00400;\
    linear1_weight_array[11][96] <= 18'h00600;\
    linear1_weight_array[11][97] <= 18'h20c00;\
    linear1_weight_array[11][98] <= 18'h00100;\
    linear1_weight_array[11][99] <= 18'h20080;\
    linear1_weight_array[11][100] <= 18'h00400;\
    linear1_weight_array[11][101] <= 18'h00600;\
    linear1_weight_array[11][102] <= 18'h20c00;\
    linear1_weight_array[11][103] <= 18'h00100;\
    linear1_weight_array[11][104] <= 18'h20080;\
    linear1_weight_array[11][105] <= 18'h00400;\
    linear1_weight_array[11][106] <= 18'h00600;\
    linear1_weight_array[11][107] <= 18'h20c00;\
    linear1_weight_array[11][108] <= 18'h00100;\
    linear1_weight_array[11][109] <= 18'h20080;\
    linear1_weight_array[11][110] <= 18'h00400;\
    linear1_weight_array[11][111] <= 18'h00600;\
    linear1_weight_array[11][112] <= 18'h20c00;\
    linear1_weight_array[11][113] <= 18'h00100;\
    linear1_weight_array[11][114] <= 18'h20080;\
    linear1_weight_array[11][115] <= 18'h00400;\
    linear1_weight_array[11][116] <= 18'h00600;\
    linear1_weight_array[11][117] <= 18'h20c00;\
    linear1_weight_array[11][118] <= 18'h00100;\
    linear1_weight_array[11][119] <= 18'h20080;\
    linear1_weight_array[11][120] <= 18'h00400;\
    linear1_weight_array[11][121] <= 18'h00600;\
    linear1_weight_array[11][122] <= 18'h20c00;\
    linear1_weight_array[11][123] <= 18'h00100;\
    linear1_weight_array[11][124] <= 18'h20080;\
    linear1_weight_array[11][125] <= 18'h00400;\
    linear1_weight_array[11][126] <= 18'h00600;\
    linear1_weight_array[11][127] <= 18'h20c00;\
    linear1_weight_array[11][128] <= 18'h00100;\
    linear1_weight_array[11][129] <= 18'h20080;\
    linear1_weight_array[11][130] <= 18'h00400;\
    linear1_weight_array[11][131] <= 18'h00600;\
    linear1_weight_array[11][132] <= 18'h20c00;\
    linear1_weight_array[11][133] <= 18'h00100;\
    linear1_weight_array[11][134] <= 18'h20080;\
    linear1_weight_array[11][135] <= 18'h00400;\
    linear1_weight_array[11][136] <= 18'h00600;\
    linear1_weight_array[11][137] <= 18'h20c00;\
    linear1_weight_array[11][138] <= 18'h00100;\
    linear1_weight_array[11][139] <= 18'h20080;\
    linear1_weight_array[11][140] <= 18'h00400;\
    linear1_weight_array[11][141] <= 18'h00600;\
    linear1_weight_array[11][142] <= 18'h20c00;\
    linear1_weight_array[11][143] <= 18'h00100;\
    linear1_weight_array[11][144] <= 18'h20080;\
    linear1_weight_array[11][145] <= 18'h00400;\
    linear1_weight_array[11][146] <= 18'h00600;\
    linear1_weight_array[11][147] <= 18'h20c00;\
    linear1_weight_array[11][148] <= 18'h00100;\
    linear1_weight_array[11][149] <= 18'h20080;\
end
*/