`define PRODUCTED \
always@(posedge clk or negedge rst_n) begin\
    if(!rst_n) begin\
		producted_1[0] <= 18'd0;\
		producted_1[1] <= 18'd0;\
		producted_1[2] <= 18'd0;\
		producted_1[3] <= 18'd0;\
		producted_1[4] <= 18'd0;\
		producted_1[5] <= 18'd0;\
		producted_1[6] <= 18'd0;\
		producted_1[7] <= 18'd0;\
		producted_1[8] <= 18'd0;\
		producted_1[9] <= 18'd0;\
		producted_1[10] <= 18'd0;\
		producted_1[11] <= 18'd0;\
		producted_1[12] <= 18'd0;\
		producted_1[13] <= 18'd0;\
		producted_1[14] <= 18'd0;\
		producted_1[15] <= 18'd0;\
		producted_1[16] <= 18'd0;\
		producted_1[17] <= 18'd0;\
		producted_1[18] <= 18'd0;\
		producted_1[19] <= 18'd0;\
		producted_1[20] <= 18'd0;\
		producted_1[21] <= 18'd0;\
		producted_1[22] <= 18'd0;\
		producted_1[23] <= 18'd0;\
		producted_1[24] <= 18'd0;\
		producted_1[25] <= 18'd0;\
		producted_1[26] <= 18'd0;\
		producted_1[27] <= 18'd0;\
		producted_1[28] <= 18'd0;\
		producted_1[29] <= 18'd0;\
		producted_1[30] <= 18'd0;\
		producted_1[31] <= 18'd0;\
		producted_1[32] <= 18'd0;\
		producted_1[33] <= 18'd0;\
		producted_1[34] <= 18'd0;\
		producted_1[35] <= 18'd0;\
		producted_1[36] <= 18'd0;\
		producted_1[37] <= 18'd0;\
		producted_1[38] <= 18'd0;\
		producted_1[39] <= 18'd0;\
		producted_1[40] <= 18'd0;\
		producted_1[41] <= 18'd0;\
		producted_1[42] <= 18'd0;\
		producted_1[43] <= 18'd0;\
		producted_1[44] <= 18'd0;\
		producted_1[45] <= 18'd0;\
		producted_1[46] <= 18'd0;\
		producted_1[47] <= 18'd0;\
		producted_1[48] <= 18'd0;\
		producted_1[49] <= 18'd0;\
		producted_1[50] <= 18'd0;\
		producted_1[51] <= 18'd0;\
		producted_1[52] <= 18'd0;\
		producted_1[53] <= 18'd0;\
		producted_1[54] <= 18'd0;\
		producted_1[55] <= 18'd0;\
		producted_1[56] <= 18'd0;\
		producted_1[57] <= 18'd0;\
		producted_1[58] <= 18'd0;\
		producted_1[59] <= 18'd0;\
		producted_1[60] <= 18'd0;\
		producted_1[61] <= 18'd0;\
		producted_1[62] <= 18'd0;\
		producted_1[63] <= 18'd0;\
		producted_1[64] <= 18'd0;\
		producted_1[65] <= 18'd0;\
		producted_1[66] <= 18'd0;\
		producted_1[67] <= 18'd0;\
		producted_1[68] <= 18'd0;\
		producted_1[69] <= 18'd0;\
		producted_1[70] <= 18'd0;\
		producted_1[71] <= 18'd0;\
		producted_1[72] <= 18'd0;\
		producted_1[73] <= 18'd0;\
		producted_1[74] <= 18'd0;\
		producted_1[75] <= 18'd0;\
		producted_1[76] <= 18'd0;\
		producted_1[77] <= 18'd0;\
		producted_1[78] <= 18'd0;\
		producted_1[79] <= 18'd0;\
		producted_1[80] <= 18'd0;\
		producted_1[81] <= 18'd0;\
		producted_1[82] <= 18'd0;\
		producted_1[83] <= 18'd0;\
		producted_1[84] <= 18'd0;\
		producted_1[85] <= 18'd0;\
		producted_1[86] <= 18'd0;\
		producted_1[87] <= 18'd0;\
		producted_1[88] <= 18'd0;\
		producted_1[89] <= 18'd0;\
		producted_1[90] <= 18'd0;\
		producted_1[91] <= 18'd0;\
		producted_1[92] <= 18'd0;\
		producted_1[93] <= 18'd0;\
		producted_1[94] <= 18'd0;\
		producted_1[95] <= 18'd0;\
		producted_1[96] <= 18'd0;\
		producted_1[97] <= 18'd0;\
		producted_1[98] <= 18'd0;\
		producted_1[99] <= 18'd0;\
		producted_1[100] <= 18'd0;\
		producted_1[101] <= 18'd0;\
		producted_1[102] <= 18'd0;\
		producted_1[103] <= 18'd0;\
		producted_1[104] <= 18'd0;\
		producted_1[105] <= 18'd0;\
		producted_1[106] <= 18'd0;\
		producted_1[107] <= 18'd0;\
		producted_1[108] <= 18'd0;\
		producted_1[109] <= 18'd0;\
		producted_1[110] <= 18'd0;\
		producted_1[111] <= 18'd0;\
    end\
    else begin\
        case(state)\
            IDLE     :;\
            INPUT    :;\
            CONV1_1_1,CONV1_2_1,CONV1_3_1,CONV1_4_1,CONV1_5_1,CONV1_6_1:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_1[0] <= in_img_array[0+cnt1][0+cnt2];\
                    producted_1[1] <= in_img_array[0+cnt1][1+cnt2];\
                    producted_1[2] <= in_img_array[0+cnt1][2+cnt2];\
                    producted_1[3] <= in_img_array[0+cnt1][3+cnt2];\
                    producted_1[4] <= in_img_array[0+cnt1][4+cnt2];\
                    producted_1[5] <= in_img_array[0+cnt1][5+cnt2];\
                    producted_1[6] <= in_img_array[0+cnt1][6+cnt2];\
                    producted_1[7] <= in_img_array[0+cnt1][7+cnt2];\
                    producted_1[8] <= in_img_array[0+cnt1][8+cnt2];\
                    producted_1[9] <= in_img_array[0+cnt1][9+cnt2];\
                    producted_1[10] <= in_img_array[0+cnt1][10+cnt2];\
                    producted_1[11] <= in_img_array[0+cnt1][11+cnt2];\
                    producted_1[12] <= in_img_array[0+cnt1][12+cnt2];\
                    producted_1[13] <= in_img_array[0+cnt1][13+cnt2];\
                    producted_1[14] <= in_img_array[0+cnt1][14+cnt2];\
                    producted_1[15] <= in_img_array[0+cnt1][15+cnt2];\
                    producted_1[16] <= in_img_array[0+cnt1][16+cnt2];\
                    producted_1[17] <= in_img_array[0+cnt1][17+cnt2];\
                    producted_1[18] <= in_img_array[0+cnt1][18+cnt2];\
                    producted_1[19] <= in_img_array[0+cnt1][19+cnt2];\
                    producted_1[20] <= in_img_array[0+cnt1][20+cnt2];\
                    producted_1[21] <= in_img_array[0+cnt1][21+cnt2];\
                    producted_1[22] <= in_img_array[0+cnt1][22+cnt2];\
                    producted_1[23] <= in_img_array[0+cnt1][23+cnt2];\
                    producted_1[24] <= in_img_array[0+cnt1][24+cnt2];\
                    producted_1[25] <= in_img_array[0+cnt1][25+cnt2];\
                    producted_1[26] <= in_img_array[0+cnt1][26+cnt2];\
                    producted_1[27] <= in_img_array[0+cnt1][27+cnt2];\
                    producted_1[28] <= in_img_array[1+cnt1][0+cnt2];\
                    producted_1[29] <= in_img_array[1+cnt1][1+cnt2];\
                    producted_1[30] <= in_img_array[1+cnt1][2+cnt2];\
                    producted_1[31] <= in_img_array[1+cnt1][3+cnt2];\
                    producted_1[32] <= in_img_array[1+cnt1][4+cnt2];\
                    producted_1[33] <= in_img_array[1+cnt1][5+cnt2];\
                    producted_1[34] <= in_img_array[1+cnt1][6+cnt2];\
                    producted_1[35] <= in_img_array[1+cnt1][7+cnt2];\
                    producted_1[36] <= in_img_array[1+cnt1][8+cnt2];\
                    producted_1[37] <= in_img_array[1+cnt1][9+cnt2];\
                    producted_1[38] <= in_img_array[1+cnt1][10+cnt2];\
                    producted_1[39] <= in_img_array[1+cnt1][11+cnt2];\
                    producted_1[40] <= in_img_array[1+cnt1][12+cnt2];\
                    producted_1[41] <= in_img_array[1+cnt1][13+cnt2];\
                    producted_1[42] <= in_img_array[1+cnt1][14+cnt2];\
                    producted_1[43] <= in_img_array[1+cnt1][15+cnt2];\
                    producted_1[44] <= in_img_array[1+cnt1][16+cnt2];\
                    producted_1[45] <= in_img_array[1+cnt1][17+cnt2];\
                    producted_1[46] <= in_img_array[1+cnt1][18+cnt2];\
                    producted_1[47] <= in_img_array[1+cnt1][19+cnt2];\
                    producted_1[48] <= in_img_array[1+cnt1][20+cnt2];\
                    producted_1[49] <= in_img_array[1+cnt1][21+cnt2];\
                    producted_1[50] <= in_img_array[1+cnt1][22+cnt2];\
                    producted_1[51] <= in_img_array[1+cnt1][23+cnt2];\
                    producted_1[52] <= in_img_array[1+cnt1][24+cnt2];\
                    producted_1[53] <= in_img_array[1+cnt1][25+cnt2];\
                    producted_1[54] <= in_img_array[1+cnt1][26+cnt2];\
                    producted_1[55] <= in_img_array[1+cnt1][27+cnt2];\
                    producted_1[56] <= in_img_array[2+cnt1][0+cnt2];\
                    producted_1[57] <= in_img_array[2+cnt1][1+cnt2];\
                    producted_1[58] <= in_img_array[2+cnt1][2+cnt2];\
                    producted_1[59] <= in_img_array[2+cnt1][3+cnt2];\
                    producted_1[60] <= in_img_array[2+cnt1][4+cnt2];\
                    producted_1[61] <= in_img_array[2+cnt1][5+cnt2];\
                    producted_1[62] <= in_img_array[2+cnt1][6+cnt2];\
                    producted_1[63] <= in_img_array[2+cnt1][7+cnt2];\
                    producted_1[64] <= in_img_array[2+cnt1][8+cnt2];\
                    producted_1[65] <= in_img_array[2+cnt1][9+cnt2];\
                    producted_1[66] <= in_img_array[2+cnt1][10+cnt2];\
                    producted_1[67] <= in_img_array[2+cnt1][11+cnt2];\
                    producted_1[68] <= in_img_array[2+cnt1][12+cnt2];\
                    producted_1[69] <= in_img_array[2+cnt1][13+cnt2];\
                    producted_1[70] <= in_img_array[2+cnt1][14+cnt2];\
                    producted_1[71] <= in_img_array[2+cnt1][15+cnt2];\
                    producted_1[72] <= in_img_array[2+cnt1][16+cnt2];\
                    producted_1[73] <= in_img_array[2+cnt1][17+cnt2];\
                    producted_1[74] <= in_img_array[2+cnt1][18+cnt2];\
                    producted_1[75] <= in_img_array[2+cnt1][19+cnt2];\
                    producted_1[76] <= in_img_array[2+cnt1][20+cnt2];\
                    producted_1[77] <= in_img_array[2+cnt1][21+cnt2];\
                    producted_1[78] <= in_img_array[2+cnt1][22+cnt2];\
                    producted_1[79] <= in_img_array[2+cnt1][23+cnt2];\
                    producted_1[80] <= in_img_array[2+cnt1][24+cnt2];\
                    producted_1[81] <= in_img_array[2+cnt1][25+cnt2];\
                    producted_1[82] <= in_img_array[2+cnt1][26+cnt2];\
                    producted_1[83] <= in_img_array[2+cnt1][27+cnt2];\
                    producted_1[84] <= in_img_array[3+cnt1][0+cnt2];\
                    producted_1[85] <= in_img_array[3+cnt1][1+cnt2];\
                    producted_1[86] <= in_img_array[3+cnt1][2+cnt2];\
                    producted_1[87] <= in_img_array[3+cnt1][3+cnt2];\
                    producted_1[88] <= in_img_array[3+cnt1][4+cnt2];\
                    producted_1[89] <= in_img_array[3+cnt1][5+cnt2];\
                    producted_1[90] <= in_img_array[3+cnt1][6+cnt2];\
                    producted_1[91] <= in_img_array[3+cnt1][7+cnt2];\
                    producted_1[92] <= in_img_array[3+cnt1][8+cnt2];\
                    producted_1[93] <= in_img_array[3+cnt1][9+cnt2];\
                    producted_1[94] <= in_img_array[3+cnt1][10+cnt2];\
                    producted_1[95] <= in_img_array[3+cnt1][11+cnt2];\
                    producted_1[96] <= in_img_array[3+cnt1][12+cnt2];\
                    producted_1[97] <= in_img_array[3+cnt1][13+cnt2];\
                    producted_1[98] <= in_img_array[3+cnt1][14+cnt2];\
                    producted_1[99] <= in_img_array[3+cnt1][15+cnt2];\
                    producted_1[100] <= in_img_array[3+cnt1][16+cnt2];\
                    producted_1[101] <= in_img_array[3+cnt1][17+cnt2];\
                    producted_1[102] <= in_img_array[3+cnt1][18+cnt2];\
                    producted_1[103] <= in_img_array[3+cnt1][19+cnt2];\
                    producted_1[104] <= in_img_array[3+cnt1][20+cnt2];\
                    producted_1[105] <= in_img_array[3+cnt1][21+cnt2];\
                    producted_1[106] <= in_img_array[3+cnt1][22+cnt2];\
                    producted_1[107] <= in_img_array[3+cnt1][23+cnt2];\
                    producted_1[108] <= in_img_array[3+cnt1][24+cnt2];\
                    producted_1[109] <= in_img_array[3+cnt1][25+cnt2];\
                    producted_1[110] <= in_img_array[3+cnt1][26+cnt2];\
                    producted_1[111] <= in_img_array[3+cnt1][27+cnt2];\
                end\
            end\
            CONV1_1_2,CONV1_2_2,CONV1_3_2,CONV1_4_2,CONV1_5_2,CONV1_6_2:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_1[0] <= in_img_array[4+cnt1][0+cnt2];\
					producted_1[1] <= in_img_array[4+cnt1][1+cnt2];\
					producted_1[2] <= in_img_array[4+cnt1][2+cnt2];\
					producted_1[3] <= in_img_array[4+cnt1][3+cnt2];\
					producted_1[4] <= in_img_array[4+cnt1][4+cnt2];\
					producted_1[5] <= in_img_array[4+cnt1][5+cnt2];\
					producted_1[6] <= in_img_array[4+cnt1][6+cnt2];\
					producted_1[7] <= in_img_array[4+cnt1][7+cnt2];\
					producted_1[8] <= in_img_array[4+cnt1][8+cnt2];\
					producted_1[9] <= in_img_array[4+cnt1][9+cnt2];\
					producted_1[10] <= in_img_array[4+cnt1][10+cnt2];\
					producted_1[11] <= in_img_array[4+cnt1][11+cnt2];\
					producted_1[12] <= in_img_array[4+cnt1][12+cnt2];\
					producted_1[13] <= in_img_array[4+cnt1][13+cnt2];\
					producted_1[14] <= in_img_array[4+cnt1][14+cnt2];\
					producted_1[15] <= in_img_array[4+cnt1][15+cnt2];\
					producted_1[16] <= in_img_array[4+cnt1][16+cnt2];\
					producted_1[17] <= in_img_array[4+cnt1][17+cnt2];\
					producted_1[18] <= in_img_array[4+cnt1][18+cnt2];\
					producted_1[19] <= in_img_array[4+cnt1][19+cnt2];\
					producted_1[20] <= in_img_array[4+cnt1][20+cnt2];\
					producted_1[21] <= in_img_array[4+cnt1][21+cnt2];\
					producted_1[22] <= in_img_array[4+cnt1][22+cnt2];\
					producted_1[23] <= in_img_array[4+cnt1][23+cnt2];\
					producted_1[24] <= in_img_array[4+cnt1][24+cnt2];\
					producted_1[25] <= in_img_array[4+cnt1][25+cnt2];\
					producted_1[26] <= in_img_array[4+cnt1][26+cnt2];\
					producted_1[27] <= in_img_array[4+cnt1][27+cnt2];\
					producted_1[28] <= in_img_array[5+cnt1][0+cnt2];\
					producted_1[29] <= in_img_array[5+cnt1][1+cnt2];\
					producted_1[30] <= in_img_array[5+cnt1][2+cnt2];\
					producted_1[31] <= in_img_array[5+cnt1][3+cnt2];\
					producted_1[32] <= in_img_array[5+cnt1][4+cnt2];\
					producted_1[33] <= in_img_array[5+cnt1][5+cnt2];\
					producted_1[34] <= in_img_array[5+cnt1][6+cnt2];\
					producted_1[35] <= in_img_array[5+cnt1][7+cnt2];\
					producted_1[36] <= in_img_array[5+cnt1][8+cnt2];\
					producted_1[37] <= in_img_array[5+cnt1][9+cnt2];\
					producted_1[38] <= in_img_array[5+cnt1][10+cnt2];\
					producted_1[39] <= in_img_array[5+cnt1][11+cnt2];\
					producted_1[40] <= in_img_array[5+cnt1][12+cnt2];\
					producted_1[41] <= in_img_array[5+cnt1][13+cnt2];\
					producted_1[42] <= in_img_array[5+cnt1][14+cnt2];\
					producted_1[43] <= in_img_array[5+cnt1][15+cnt2];\
					producted_1[44] <= in_img_array[5+cnt1][16+cnt2];\
					producted_1[45] <= in_img_array[5+cnt1][17+cnt2];\
					producted_1[46] <= in_img_array[5+cnt1][18+cnt2];\
					producted_1[47] <= in_img_array[5+cnt1][19+cnt2];\
					producted_1[48] <= in_img_array[5+cnt1][20+cnt2];\
					producted_1[49] <= in_img_array[5+cnt1][21+cnt2];\
					producted_1[50] <= in_img_array[5+cnt1][22+cnt2];\
					producted_1[51] <= in_img_array[5+cnt1][23+cnt2];\
					producted_1[52] <= in_img_array[5+cnt1][24+cnt2];\
					producted_1[53] <= in_img_array[5+cnt1][25+cnt2];\
					producted_1[54] <= in_img_array[5+cnt1][26+cnt2];\
					producted_1[55] <= in_img_array[5+cnt1][27+cnt2];\
					producted_1[56] <= in_img_array[6+cnt1][0+cnt2];\
					producted_1[57] <= in_img_array[6+cnt1][1+cnt2];\
					producted_1[58] <= in_img_array[6+cnt1][2+cnt2];\
					producted_1[59] <= in_img_array[6+cnt1][3+cnt2];\
					producted_1[60] <= in_img_array[6+cnt1][4+cnt2];\
					producted_1[61] <= in_img_array[6+cnt1][5+cnt2];\
					producted_1[62] <= in_img_array[6+cnt1][6+cnt2];\
					producted_1[63] <= in_img_array[6+cnt1][7+cnt2];\
					producted_1[64] <= in_img_array[6+cnt1][8+cnt2];\
					producted_1[65] <= in_img_array[6+cnt1][9+cnt2];\
					producted_1[66] <= in_img_array[6+cnt1][10+cnt2];\
					producted_1[67] <= in_img_array[6+cnt1][11+cnt2];\
					producted_1[68] <= in_img_array[6+cnt1][12+cnt2];\
					producted_1[69] <= in_img_array[6+cnt1][13+cnt2];\
					producted_1[70] <= in_img_array[6+cnt1][14+cnt2];\
					producted_1[71] <= in_img_array[6+cnt1][15+cnt2];\
					producted_1[72] <= in_img_array[6+cnt1][16+cnt2];\
					producted_1[73] <= in_img_array[6+cnt1][17+cnt2];\
					producted_1[74] <= in_img_array[6+cnt1][18+cnt2];\
					producted_1[75] <= in_img_array[6+cnt1][19+cnt2];\
					producted_1[76] <= in_img_array[6+cnt1][20+cnt2];\
					producted_1[77] <= in_img_array[6+cnt1][21+cnt2];\
					producted_1[78] <= in_img_array[6+cnt1][22+cnt2];\
					producted_1[79] <= in_img_array[6+cnt1][23+cnt2];\
					producted_1[80] <= in_img_array[6+cnt1][24+cnt2];\
					producted_1[81] <= in_img_array[6+cnt1][25+cnt2];\
					producted_1[82] <= in_img_array[6+cnt1][26+cnt2];\
					producted_1[83] <= in_img_array[6+cnt1][27+cnt2];\
					producted_1[84] <= in_img_array[7+cnt1][0+cnt2];\
					producted_1[85] <= in_img_array[7+cnt1][1+cnt2];\
					producted_1[86] <= in_img_array[7+cnt1][2+cnt2];\
					producted_1[87] <= in_img_array[7+cnt1][3+cnt2];\
					producted_1[88] <= in_img_array[7+cnt1][4+cnt2];\
					producted_1[89] <= in_img_array[7+cnt1][5+cnt2];\
					producted_1[90] <= in_img_array[7+cnt1][6+cnt2];\
					producted_1[91] <= in_img_array[7+cnt1][7+cnt2];\
					producted_1[92] <= in_img_array[7+cnt1][8+cnt2];\
					producted_1[93] <= in_img_array[7+cnt1][9+cnt2];\
					producted_1[94] <= in_img_array[7+cnt1][10+cnt2];\
					producted_1[95] <= in_img_array[7+cnt1][11+cnt2];\
					producted_1[96] <= in_img_array[7+cnt1][12+cnt2];\
					producted_1[97] <= in_img_array[7+cnt1][13+cnt2];\
					producted_1[98] <= in_img_array[7+cnt1][14+cnt2];\
					producted_1[99] <= in_img_array[7+cnt1][15+cnt2];\
					producted_1[100] <= in_img_array[7+cnt1][16+cnt2];\
					producted_1[101] <= in_img_array[7+cnt1][17+cnt2];\
					producted_1[102] <= in_img_array[7+cnt1][18+cnt2];\
					producted_1[103] <= in_img_array[7+cnt1][19+cnt2];\
					producted_1[104] <= in_img_array[7+cnt1][20+cnt2];\
					producted_1[105] <= in_img_array[7+cnt1][21+cnt2];\
					producted_1[106] <= in_img_array[7+cnt1][22+cnt2];\
					producted_1[107] <= in_img_array[7+cnt1][23+cnt2];\
					producted_1[108] <= in_img_array[7+cnt1][24+cnt2];\
					producted_1[109] <= in_img_array[7+cnt1][25+cnt2];\
					producted_1[110] <= in_img_array[7+cnt1][26+cnt2];\
					producted_1[111] <= in_img_array[7+cnt1][27+cnt2];\
                end\
            end\
            CONV1_1_3,CONV1_2_3,CONV1_3_3,CONV1_4_3,CONV1_5_3,CONV1_6_3:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_1[0] <= in_img_array[8+cnt1][0+cnt2];\
					producted_1[1] <= in_img_array[8+cnt1][1+cnt2];\
					producted_1[2] <= in_img_array[8+cnt1][2+cnt2];\
					producted_1[3] <= in_img_array[8+cnt1][3+cnt2];\
					producted_1[4] <= in_img_array[8+cnt1][4+cnt2];\
					producted_1[5] <= in_img_array[8+cnt1][5+cnt2];\
					producted_1[6] <= in_img_array[8+cnt1][6+cnt2];\
					producted_1[7] <= in_img_array[8+cnt1][7+cnt2];\
					producted_1[8] <= in_img_array[8+cnt1][8+cnt2];\
					producted_1[9] <= in_img_array[8+cnt1][9+cnt2];\
					producted_1[10] <= in_img_array[8+cnt1][10+cnt2];\
					producted_1[11] <= in_img_array[8+cnt1][11+cnt2];\
					producted_1[12] <= in_img_array[8+cnt1][12+cnt2];\
					producted_1[13] <= in_img_array[8+cnt1][13+cnt2];\
					producted_1[14] <= in_img_array[8+cnt1][14+cnt2];\
					producted_1[15] <= in_img_array[8+cnt1][15+cnt2];\
					producted_1[16] <= in_img_array[8+cnt1][16+cnt2];\
					producted_1[17] <= in_img_array[8+cnt1][17+cnt2];\
					producted_1[18] <= in_img_array[8+cnt1][18+cnt2];\
					producted_1[19] <= in_img_array[8+cnt1][19+cnt2];\
					producted_1[20] <= in_img_array[8+cnt1][20+cnt2];\
					producted_1[21] <= in_img_array[8+cnt1][21+cnt2];\
					producted_1[22] <= in_img_array[8+cnt1][22+cnt2];\
					producted_1[23] <= in_img_array[8+cnt1][23+cnt2];\
					producted_1[24] <= in_img_array[8+cnt1][24+cnt2];\
					producted_1[25] <= in_img_array[8+cnt1][25+cnt2];\
					producted_1[26] <= in_img_array[8+cnt1][26+cnt2];\
					producted_1[27] <= in_img_array[8+cnt1][27+cnt2];\
					producted_1[28] <= in_img_array[9+cnt1][0+cnt2];\
					producted_1[29] <= in_img_array[9+cnt1][1+cnt2];\
					producted_1[30] <= in_img_array[9+cnt1][2+cnt2];\
					producted_1[31] <= in_img_array[9+cnt1][3+cnt2];\
					producted_1[32] <= in_img_array[9+cnt1][4+cnt2];\
					producted_1[33] <= in_img_array[9+cnt1][5+cnt2];\
					producted_1[34] <= in_img_array[9+cnt1][6+cnt2];\
					producted_1[35] <= in_img_array[9+cnt1][7+cnt2];\
					producted_1[36] <= in_img_array[9+cnt1][8+cnt2];\
					producted_1[37] <= in_img_array[9+cnt1][9+cnt2];\
					producted_1[38] <= in_img_array[9+cnt1][10+cnt2];\
					producted_1[39] <= in_img_array[9+cnt1][11+cnt2];\
					producted_1[40] <= in_img_array[9+cnt1][12+cnt2];\
					producted_1[41] <= in_img_array[9+cnt1][13+cnt2];\
					producted_1[42] <= in_img_array[9+cnt1][14+cnt2];\
					producted_1[43] <= in_img_array[9+cnt1][15+cnt2];\
					producted_1[44] <= in_img_array[9+cnt1][16+cnt2];\
					producted_1[45] <= in_img_array[9+cnt1][17+cnt2];\
					producted_1[46] <= in_img_array[9+cnt1][18+cnt2];\
					producted_1[47] <= in_img_array[9+cnt1][19+cnt2];\
					producted_1[48] <= in_img_array[9+cnt1][20+cnt2];\
					producted_1[49] <= in_img_array[9+cnt1][21+cnt2];\
					producted_1[50] <= in_img_array[9+cnt1][22+cnt2];\
					producted_1[51] <= in_img_array[9+cnt1][23+cnt2];\
					producted_1[52] <= in_img_array[9+cnt1][24+cnt2];\
					producted_1[53] <= in_img_array[9+cnt1][25+cnt2];\
					producted_1[54] <= in_img_array[9+cnt1][26+cnt2];\
					producted_1[55] <= in_img_array[9+cnt1][27+cnt2];\
					producted_1[56] <= in_img_array[10+cnt1][0+cnt2];\
					producted_1[57] <= in_img_array[10+cnt1][1+cnt2];\
					producted_1[58] <= in_img_array[10+cnt1][2+cnt2];\
					producted_1[59] <= in_img_array[10+cnt1][3+cnt2];\
					producted_1[60] <= in_img_array[10+cnt1][4+cnt2];\
					producted_1[61] <= in_img_array[10+cnt1][5+cnt2];\
					producted_1[62] <= in_img_array[10+cnt1][6+cnt2];\
					producted_1[63] <= in_img_array[10+cnt1][7+cnt2];\
					producted_1[64] <= in_img_array[10+cnt1][8+cnt2];\
					producted_1[65] <= in_img_array[10+cnt1][9+cnt2];\
					producted_1[66] <= in_img_array[10+cnt1][10+cnt2];\
					producted_1[67] <= in_img_array[10+cnt1][11+cnt2];\
					producted_1[68] <= in_img_array[10+cnt1][12+cnt2];\
					producted_1[69] <= in_img_array[10+cnt1][13+cnt2];\
					producted_1[70] <= in_img_array[10+cnt1][14+cnt2];\
					producted_1[71] <= in_img_array[10+cnt1][15+cnt2];\
					producted_1[72] <= in_img_array[10+cnt1][16+cnt2];\
					producted_1[73] <= in_img_array[10+cnt1][17+cnt2];\
					producted_1[74] <= in_img_array[10+cnt1][18+cnt2];\
					producted_1[75] <= in_img_array[10+cnt1][19+cnt2];\
					producted_1[76] <= in_img_array[10+cnt1][20+cnt2];\
					producted_1[77] <= in_img_array[10+cnt1][21+cnt2];\
					producted_1[78] <= in_img_array[10+cnt1][22+cnt2];\
					producted_1[79] <= in_img_array[10+cnt1][23+cnt2];\
					producted_1[80] <= in_img_array[10+cnt1][24+cnt2];\
					producted_1[81] <= in_img_array[10+cnt1][25+cnt2];\
					producted_1[82] <= in_img_array[10+cnt1][26+cnt2];\
					producted_1[83] <= in_img_array[10+cnt1][27+cnt2];\
					producted_1[84] <= in_img_array[11+cnt1][0+cnt2];\
					producted_1[85] <= in_img_array[11+cnt1][1+cnt2];\
					producted_1[86] <= in_img_array[11+cnt1][2+cnt2];\
					producted_1[87] <= in_img_array[11+cnt1][3+cnt2];\
					producted_1[88] <= in_img_array[11+cnt1][4+cnt2];\
					producted_1[89] <= in_img_array[11+cnt1][5+cnt2];\
					producted_1[90] <= in_img_array[11+cnt1][6+cnt2];\
					producted_1[91] <= in_img_array[11+cnt1][7+cnt2];\
					producted_1[92] <= in_img_array[11+cnt1][8+cnt2];\
					producted_1[93] <= in_img_array[11+cnt1][9+cnt2];\
					producted_1[94] <= in_img_array[11+cnt1][10+cnt2];\
					producted_1[95] <= in_img_array[11+cnt1][11+cnt2];\
					producted_1[96] <= in_img_array[11+cnt1][12+cnt2];\
					producted_1[97] <= in_img_array[11+cnt1][13+cnt2];\
					producted_1[98] <= in_img_array[11+cnt1][14+cnt2];\
					producted_1[99] <= in_img_array[11+cnt1][15+cnt2];\
					producted_1[100] <= in_img_array[11+cnt1][16+cnt2];\
					producted_1[101] <= in_img_array[11+cnt1][17+cnt2];\
					producted_1[102] <= in_img_array[11+cnt1][18+cnt2];\
					producted_1[103] <= in_img_array[11+cnt1][19+cnt2];\
					producted_1[104] <= in_img_array[11+cnt1][20+cnt2];\
					producted_1[105] <= in_img_array[11+cnt1][21+cnt2];\
					producted_1[106] <= in_img_array[11+cnt1][22+cnt2];\
					producted_1[107] <= in_img_array[11+cnt1][23+cnt2];\
					producted_1[108] <= in_img_array[11+cnt1][24+cnt2];\
					producted_1[109] <= in_img_array[11+cnt1][25+cnt2];\
					producted_1[110] <= in_img_array[11+cnt1][26+cnt2];\
					producted_1[111] <= in_img_array[11+cnt1][27+cnt2];\
                end\
            end\
            CONV1_1_4,CONV1_2_4,CONV1_3_4,CONV1_4_4,CONV1_5_4,CONV1_6_4:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_1[0] <= in_img_array[12+cnt1][0+cnt2];\
					producted_1[1] <= in_img_array[12+cnt1][1+cnt2];\
					producted_1[2] <= in_img_array[12+cnt1][2+cnt2];\
					producted_1[3] <= in_img_array[12+cnt1][3+cnt2];\
					producted_1[4] <= in_img_array[12+cnt1][4+cnt2];\
					producted_1[5] <= in_img_array[12+cnt1][5+cnt2];\
					producted_1[6] <= in_img_array[12+cnt1][6+cnt2];\
					producted_1[7] <= in_img_array[12+cnt1][7+cnt2];\
					producted_1[8] <= in_img_array[12+cnt1][8+cnt2];\
					producted_1[9] <= in_img_array[12+cnt1][9+cnt2];\
					producted_1[10] <= in_img_array[12+cnt1][10+cnt2];\
					producted_1[11] <= in_img_array[12+cnt1][11+cnt2];\
					producted_1[12] <= in_img_array[12+cnt1][12+cnt2];\
					producted_1[13] <= in_img_array[12+cnt1][13+cnt2];\
					producted_1[14] <= in_img_array[12+cnt1][14+cnt2];\
					producted_1[15] <= in_img_array[12+cnt1][15+cnt2];\
					producted_1[16] <= in_img_array[12+cnt1][16+cnt2];\
					producted_1[17] <= in_img_array[12+cnt1][17+cnt2];\
					producted_1[18] <= in_img_array[12+cnt1][18+cnt2];\
					producted_1[19] <= in_img_array[12+cnt1][19+cnt2];\
					producted_1[20] <= in_img_array[12+cnt1][20+cnt2];\
					producted_1[21] <= in_img_array[12+cnt1][21+cnt2];\
					producted_1[22] <= in_img_array[12+cnt1][22+cnt2];\
					producted_1[23] <= in_img_array[12+cnt1][23+cnt2];\
					producted_1[24] <= in_img_array[12+cnt1][24+cnt2];\
					producted_1[25] <= in_img_array[12+cnt1][25+cnt2];\
					producted_1[26] <= in_img_array[12+cnt1][26+cnt2];\
					producted_1[27] <= in_img_array[12+cnt1][27+cnt2];\
					producted_1[28] <= in_img_array[13+cnt1][0+cnt2];\
					producted_1[29] <= in_img_array[13+cnt1][1+cnt2];\
					producted_1[30] <= in_img_array[13+cnt1][2+cnt2];\
					producted_1[31] <= in_img_array[13+cnt1][3+cnt2];\
					producted_1[32] <= in_img_array[13+cnt1][4+cnt2];\
					producted_1[33] <= in_img_array[13+cnt1][5+cnt2];\
					producted_1[34] <= in_img_array[13+cnt1][6+cnt2];\
					producted_1[35] <= in_img_array[13+cnt1][7+cnt2];\
					producted_1[36] <= in_img_array[13+cnt1][8+cnt2];\
					producted_1[37] <= in_img_array[13+cnt1][9+cnt2];\
					producted_1[38] <= in_img_array[13+cnt1][10+cnt2];\
					producted_1[39] <= in_img_array[13+cnt1][11+cnt2];\
					producted_1[40] <= in_img_array[13+cnt1][12+cnt2];\
					producted_1[41] <= in_img_array[13+cnt1][13+cnt2];\
					producted_1[42] <= in_img_array[13+cnt1][14+cnt2];\
					producted_1[43] <= in_img_array[13+cnt1][15+cnt2];\
					producted_1[44] <= in_img_array[13+cnt1][16+cnt2];\
					producted_1[45] <= in_img_array[13+cnt1][17+cnt2];\
					producted_1[46] <= in_img_array[13+cnt1][18+cnt2];\
					producted_1[47] <= in_img_array[13+cnt1][19+cnt2];\
					producted_1[48] <= in_img_array[13+cnt1][20+cnt2];\
					producted_1[49] <= in_img_array[13+cnt1][21+cnt2];\
					producted_1[50] <= in_img_array[13+cnt1][22+cnt2];\
					producted_1[51] <= in_img_array[13+cnt1][23+cnt2];\
					producted_1[52] <= in_img_array[13+cnt1][24+cnt2];\
					producted_1[53] <= in_img_array[13+cnt1][25+cnt2];\
					producted_1[54] <= in_img_array[13+cnt1][26+cnt2];\
					producted_1[55] <= in_img_array[13+cnt1][27+cnt2];\
					producted_1[56] <= in_img_array[14+cnt1][0+cnt2];\
					producted_1[57] <= in_img_array[14+cnt1][1+cnt2];\
					producted_1[58] <= in_img_array[14+cnt1][2+cnt2];\
					producted_1[59] <= in_img_array[14+cnt1][3+cnt2];\
					producted_1[60] <= in_img_array[14+cnt1][4+cnt2];\
					producted_1[61] <= in_img_array[14+cnt1][5+cnt2];\
					producted_1[62] <= in_img_array[14+cnt1][6+cnt2];\
					producted_1[63] <= in_img_array[14+cnt1][7+cnt2];\
					producted_1[64] <= in_img_array[14+cnt1][8+cnt2];\
					producted_1[65] <= in_img_array[14+cnt1][9+cnt2];\
					producted_1[66] <= in_img_array[14+cnt1][10+cnt2];\
					producted_1[67] <= in_img_array[14+cnt1][11+cnt2];\
					producted_1[68] <= in_img_array[14+cnt1][12+cnt2];\
					producted_1[69] <= in_img_array[14+cnt1][13+cnt2];\
					producted_1[70] <= in_img_array[14+cnt1][14+cnt2];\
					producted_1[71] <= in_img_array[14+cnt1][15+cnt2];\
					producted_1[72] <= in_img_array[14+cnt1][16+cnt2];\
					producted_1[73] <= in_img_array[14+cnt1][17+cnt2];\
					producted_1[74] <= in_img_array[14+cnt1][18+cnt2];\
					producted_1[75] <= in_img_array[14+cnt1][19+cnt2];\
					producted_1[76] <= in_img_array[14+cnt1][20+cnt2];\
					producted_1[77] <= in_img_array[14+cnt1][21+cnt2];\
					producted_1[78] <= in_img_array[14+cnt1][22+cnt2];\
					producted_1[79] <= in_img_array[14+cnt1][23+cnt2];\
					producted_1[80] <= in_img_array[14+cnt1][24+cnt2];\
					producted_1[81] <= in_img_array[14+cnt1][25+cnt2];\
					producted_1[82] <= in_img_array[14+cnt1][26+cnt2];\
					producted_1[83] <= in_img_array[14+cnt1][27+cnt2];\
					producted_1[84] <= in_img_array[15+cnt1][0+cnt2];\
					producted_1[85] <= in_img_array[15+cnt1][1+cnt2];\
					producted_1[86] <= in_img_array[15+cnt1][2+cnt2];\
					producted_1[87] <= in_img_array[15+cnt1][3+cnt2];\
					producted_1[88] <= in_img_array[15+cnt1][4+cnt2];\
					producted_1[89] <= in_img_array[15+cnt1][5+cnt2];\
					producted_1[90] <= in_img_array[15+cnt1][6+cnt2];\
					producted_1[91] <= in_img_array[15+cnt1][7+cnt2];\
					producted_1[92] <= in_img_array[15+cnt1][8+cnt2];\
					producted_1[93] <= in_img_array[15+cnt1][9+cnt2];\
					producted_1[94] <= in_img_array[15+cnt1][10+cnt2];\
					producted_1[95] <= in_img_array[15+cnt1][11+cnt2];\
					producted_1[96] <= in_img_array[15+cnt1][12+cnt2];\
					producted_1[97] <= in_img_array[15+cnt1][13+cnt2];\
					producted_1[98] <= in_img_array[15+cnt1][14+cnt2];\
					producted_1[99] <= in_img_array[15+cnt1][15+cnt2];\
					producted_1[100] <= in_img_array[15+cnt1][16+cnt2];\
					producted_1[101] <= in_img_array[15+cnt1][17+cnt2];\
					producted_1[102] <= in_img_array[15+cnt1][18+cnt2];\
					producted_1[103] <= in_img_array[15+cnt1][19+cnt2];\
					producted_1[104] <= in_img_array[15+cnt1][20+cnt2];\
					producted_1[105] <= in_img_array[15+cnt1][21+cnt2];\
					producted_1[106] <= in_img_array[15+cnt1][22+cnt2];\
					producted_1[107] <= in_img_array[15+cnt1][23+cnt2];\
					producted_1[108] <= in_img_array[15+cnt1][24+cnt2];\
					producted_1[109] <= in_img_array[15+cnt1][25+cnt2];\
					producted_1[110] <= in_img_array[15+cnt1][26+cnt2];\
					producted_1[111] <= in_img_array[15+cnt1][27+cnt2];\
                end\
            end\
            CONV1_1_5,CONV1_2_5,CONV1_3_5,CONV1_4_5,CONV1_5_5,CONV1_6_5:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_1[0] <= in_img_array[16+cnt1][0+cnt2];\
					producted_1[1] <= in_img_array[16+cnt1][1+cnt2];\
					producted_1[2] <= in_img_array[16+cnt1][2+cnt2];\
					producted_1[3] <= in_img_array[16+cnt1][3+cnt2];\
					producted_1[4] <= in_img_array[16+cnt1][4+cnt2];\
					producted_1[5] <= in_img_array[16+cnt1][5+cnt2];\
					producted_1[6] <= in_img_array[16+cnt1][6+cnt2];\
					producted_1[7] <= in_img_array[16+cnt1][7+cnt2];\
					producted_1[8] <= in_img_array[16+cnt1][8+cnt2];\
					producted_1[9] <= in_img_array[16+cnt1][9+cnt2];\
					producted_1[10] <= in_img_array[16+cnt1][10+cnt2];\
					producted_1[11] <= in_img_array[16+cnt1][11+cnt2];\
					producted_1[12] <= in_img_array[16+cnt1][12+cnt2];\
					producted_1[13] <= in_img_array[16+cnt1][13+cnt2];\
					producted_1[14] <= in_img_array[16+cnt1][14+cnt2];\
					producted_1[15] <= in_img_array[16+cnt1][15+cnt2];\
					producted_1[16] <= in_img_array[16+cnt1][16+cnt2];\
					producted_1[17] <= in_img_array[16+cnt1][17+cnt2];\
					producted_1[18] <= in_img_array[16+cnt1][18+cnt2];\
					producted_1[19] <= in_img_array[16+cnt1][19+cnt2];\
					producted_1[20] <= in_img_array[16+cnt1][20+cnt2];\
					producted_1[21] <= in_img_array[16+cnt1][21+cnt2];\
					producted_1[22] <= in_img_array[16+cnt1][22+cnt2];\
					producted_1[23] <= in_img_array[16+cnt1][23+cnt2];\
					producted_1[24] <= in_img_array[16+cnt1][24+cnt2];\
					producted_1[25] <= in_img_array[16+cnt1][25+cnt2];\
					producted_1[26] <= in_img_array[16+cnt1][26+cnt2];\
					producted_1[27] <= in_img_array[16+cnt1][27+cnt2];\
					producted_1[28] <= in_img_array[17+cnt1][0+cnt2];\
					producted_1[29] <= in_img_array[17+cnt1][1+cnt2];\
					producted_1[30] <= in_img_array[17+cnt1][2+cnt2];\
					producted_1[31] <= in_img_array[17+cnt1][3+cnt2];\
					producted_1[32] <= in_img_array[17+cnt1][4+cnt2];\
					producted_1[33] <= in_img_array[17+cnt1][5+cnt2];\
					producted_1[34] <= in_img_array[17+cnt1][6+cnt2];\
					producted_1[35] <= in_img_array[17+cnt1][7+cnt2];\
					producted_1[36] <= in_img_array[17+cnt1][8+cnt2];\
					producted_1[37] <= in_img_array[17+cnt1][9+cnt2];\
					producted_1[38] <= in_img_array[17+cnt1][10+cnt2];\
					producted_1[39] <= in_img_array[17+cnt1][11+cnt2];\
					producted_1[40] <= in_img_array[17+cnt1][12+cnt2];\
					producted_1[41] <= in_img_array[17+cnt1][13+cnt2];\
					producted_1[42] <= in_img_array[17+cnt1][14+cnt2];\
					producted_1[43] <= in_img_array[17+cnt1][15+cnt2];\
					producted_1[44] <= in_img_array[17+cnt1][16+cnt2];\
					producted_1[45] <= in_img_array[17+cnt1][17+cnt2];\
					producted_1[46] <= in_img_array[17+cnt1][18+cnt2];\
					producted_1[47] <= in_img_array[17+cnt1][19+cnt2];\
					producted_1[48] <= in_img_array[17+cnt1][20+cnt2];\
					producted_1[49] <= in_img_array[17+cnt1][21+cnt2];\
					producted_1[50] <= in_img_array[17+cnt1][22+cnt2];\
					producted_1[51] <= in_img_array[17+cnt1][23+cnt2];\
					producted_1[52] <= in_img_array[17+cnt1][24+cnt2];\
					producted_1[53] <= in_img_array[17+cnt1][25+cnt2];\
					producted_1[54] <= in_img_array[17+cnt1][26+cnt2];\
					producted_1[55] <= in_img_array[17+cnt1][27+cnt2];\
					producted_1[56] <= in_img_array[18+cnt1][0+cnt2];\
					producted_1[57] <= in_img_array[18+cnt1][1+cnt2];\
					producted_1[58] <= in_img_array[18+cnt1][2+cnt2];\
					producted_1[59] <= in_img_array[18+cnt1][3+cnt2];\
					producted_1[60] <= in_img_array[18+cnt1][4+cnt2];\
					producted_1[61] <= in_img_array[18+cnt1][5+cnt2];\
					producted_1[62] <= in_img_array[18+cnt1][6+cnt2];\
					producted_1[63] <= in_img_array[18+cnt1][7+cnt2];\
					producted_1[64] <= in_img_array[18+cnt1][8+cnt2];\
					producted_1[65] <= in_img_array[18+cnt1][9+cnt2];\
					producted_1[66] <= in_img_array[18+cnt1][10+cnt2];\
					producted_1[67] <= in_img_array[18+cnt1][11+cnt2];\
					producted_1[68] <= in_img_array[18+cnt1][12+cnt2];\
					producted_1[69] <= in_img_array[18+cnt1][13+cnt2];\
					producted_1[70] <= in_img_array[18+cnt1][14+cnt2];\
					producted_1[71] <= in_img_array[18+cnt1][15+cnt2];\
					producted_1[72] <= in_img_array[18+cnt1][16+cnt2];\
					producted_1[73] <= in_img_array[18+cnt1][17+cnt2];\
					producted_1[74] <= in_img_array[18+cnt1][18+cnt2];\
					producted_1[75] <= in_img_array[18+cnt1][19+cnt2];\
					producted_1[76] <= in_img_array[18+cnt1][20+cnt2];\
					producted_1[77] <= in_img_array[18+cnt1][21+cnt2];\
					producted_1[78] <= in_img_array[18+cnt1][22+cnt2];\
					producted_1[79] <= in_img_array[18+cnt1][23+cnt2];\
					producted_1[80] <= in_img_array[18+cnt1][24+cnt2];\
					producted_1[81] <= in_img_array[18+cnt1][25+cnt2];\
					producted_1[82] <= in_img_array[18+cnt1][26+cnt2];\
					producted_1[83] <= in_img_array[18+cnt1][27+cnt2];\
					producted_1[84] <= in_img_array[19+cnt1][0+cnt2];\
					producted_1[85] <= in_img_array[19+cnt1][1+cnt2];\
					producted_1[86] <= in_img_array[19+cnt1][2+cnt2];\
					producted_1[87] <= in_img_array[19+cnt1][3+cnt2];\
					producted_1[88] <= in_img_array[19+cnt1][4+cnt2];\
					producted_1[89] <= in_img_array[19+cnt1][5+cnt2];\
					producted_1[90] <= in_img_array[19+cnt1][6+cnt2];\
					producted_1[91] <= in_img_array[19+cnt1][7+cnt2];\
					producted_1[92] <= in_img_array[19+cnt1][8+cnt2];\
					producted_1[93] <= in_img_array[19+cnt1][9+cnt2];\
					producted_1[94] <= in_img_array[19+cnt1][10+cnt2];\
					producted_1[95] <= in_img_array[19+cnt1][11+cnt2];\
					producted_1[96] <= in_img_array[19+cnt1][12+cnt2];\
					producted_1[97] <= in_img_array[19+cnt1][13+cnt2];\
					producted_1[98] <= in_img_array[19+cnt1][14+cnt2];\
					producted_1[99] <= in_img_array[19+cnt1][15+cnt2];\
					producted_1[100] <= in_img_array[19+cnt1][16+cnt2];\
					producted_1[101] <= in_img_array[19+cnt1][17+cnt2];\
					producted_1[102] <= in_img_array[19+cnt1][18+cnt2];\
					producted_1[103] <= in_img_array[19+cnt1][19+cnt2];\
					producted_1[104] <= in_img_array[19+cnt1][20+cnt2];\
					producted_1[105] <= in_img_array[19+cnt1][21+cnt2];\
					producted_1[106] <= in_img_array[19+cnt1][22+cnt2];\
					producted_1[107] <= in_img_array[19+cnt1][23+cnt2];\
					producted_1[108] <= in_img_array[19+cnt1][24+cnt2];\
					producted_1[109] <= in_img_array[19+cnt1][25+cnt2];\
					producted_1[110] <= in_img_array[19+cnt1][26+cnt2];\
					producted_1[111] <= in_img_array[19+cnt1][27+cnt2];\
                end\
            end\
            CONV1_1_6,CONV1_2_6,CONV1_3_6,CONV1_4_6,CONV1_5_6,CONV1_6_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_1[0] <= in_img_array[20+cnt1][0+cnt2];\
					producted_1[1] <= in_img_array[20+cnt1][1+cnt2];\
					producted_1[2] <= in_img_array[20+cnt1][2+cnt2];\
					producted_1[3] <= in_img_array[20+cnt1][3+cnt2];\
					producted_1[4] <= in_img_array[20+cnt1][4+cnt2];\
					producted_1[5] <= in_img_array[20+cnt1][5+cnt2];\
					producted_1[6] <= in_img_array[20+cnt1][6+cnt2];\
					producted_1[7] <= in_img_array[20+cnt1][7+cnt2];\
					producted_1[8] <= in_img_array[20+cnt1][8+cnt2];\
					producted_1[9] <= in_img_array[20+cnt1][9+cnt2];\
					producted_1[10] <= in_img_array[20+cnt1][10+cnt2];\
					producted_1[11] <= in_img_array[20+cnt1][11+cnt2];\
					producted_1[12] <= in_img_array[20+cnt1][12+cnt2];\
					producted_1[13] <= in_img_array[20+cnt1][13+cnt2];\
					producted_1[14] <= in_img_array[20+cnt1][14+cnt2];\
					producted_1[15] <= in_img_array[20+cnt1][15+cnt2];\
					producted_1[16] <= in_img_array[20+cnt1][16+cnt2];\
					producted_1[17] <= in_img_array[20+cnt1][17+cnt2];\
					producted_1[18] <= in_img_array[20+cnt1][18+cnt2];\
					producted_1[19] <= in_img_array[20+cnt1][19+cnt2];\
					producted_1[20] <= in_img_array[20+cnt1][20+cnt2];\
					producted_1[21] <= in_img_array[20+cnt1][21+cnt2];\
					producted_1[22] <= in_img_array[20+cnt1][22+cnt2];\
					producted_1[23] <= in_img_array[20+cnt1][23+cnt2];\
					producted_1[24] <= in_img_array[20+cnt1][24+cnt2];\
					producted_1[25] <= in_img_array[20+cnt1][25+cnt2];\
					producted_1[26] <= in_img_array[20+cnt1][26+cnt2];\
					producted_1[27] <= in_img_array[20+cnt1][27+cnt2];\
					producted_1[28] <= in_img_array[21+cnt1][0+cnt2];\
					producted_1[29] <= in_img_array[21+cnt1][1+cnt2];\
					producted_1[30] <= in_img_array[21+cnt1][2+cnt2];\
					producted_1[31] <= in_img_array[21+cnt1][3+cnt2];\
					producted_1[32] <= in_img_array[21+cnt1][4+cnt2];\
					producted_1[33] <= in_img_array[21+cnt1][5+cnt2];\
					producted_1[34] <= in_img_array[21+cnt1][6+cnt2];\
					producted_1[35] <= in_img_array[21+cnt1][7+cnt2];\
					producted_1[36] <= in_img_array[21+cnt1][8+cnt2];\
					producted_1[37] <= in_img_array[21+cnt1][9+cnt2];\
					producted_1[38] <= in_img_array[21+cnt1][10+cnt2];\
					producted_1[39] <= in_img_array[21+cnt1][11+cnt2];\
					producted_1[40] <= in_img_array[21+cnt1][12+cnt2];\
					producted_1[41] <= in_img_array[21+cnt1][13+cnt2];\
					producted_1[42] <= in_img_array[21+cnt1][14+cnt2];\
					producted_1[43] <= in_img_array[21+cnt1][15+cnt2];\
					producted_1[44] <= in_img_array[21+cnt1][16+cnt2];\
					producted_1[45] <= in_img_array[21+cnt1][17+cnt2];\
					producted_1[46] <= in_img_array[21+cnt1][18+cnt2];\
					producted_1[47] <= in_img_array[21+cnt1][19+cnt2];\
					producted_1[48] <= in_img_array[21+cnt1][20+cnt2];\
					producted_1[49] <= in_img_array[21+cnt1][21+cnt2];\
					producted_1[50] <= in_img_array[21+cnt1][22+cnt2];\
					producted_1[51] <= in_img_array[21+cnt1][23+cnt2];\
					producted_1[52] <= in_img_array[21+cnt1][24+cnt2];\
					producted_1[53] <= in_img_array[21+cnt1][25+cnt2];\
					producted_1[54] <= in_img_array[21+cnt1][26+cnt2];\
					producted_1[55] <= in_img_array[21+cnt1][27+cnt2];\
					producted_1[56] <= in_img_array[22+cnt1][0+cnt2];\
					producted_1[57] <= in_img_array[22+cnt1][1+cnt2];\
					producted_1[58] <= in_img_array[22+cnt1][2+cnt2];\
					producted_1[59] <= in_img_array[22+cnt1][3+cnt2];\
					producted_1[60] <= in_img_array[22+cnt1][4+cnt2];\
					producted_1[61] <= in_img_array[22+cnt1][5+cnt2];\
					producted_1[62] <= in_img_array[22+cnt1][6+cnt2];\
					producted_1[63] <= in_img_array[22+cnt1][7+cnt2];\
					producted_1[64] <= in_img_array[22+cnt1][8+cnt2];\
					producted_1[65] <= in_img_array[22+cnt1][9+cnt2];\
					producted_1[66] <= in_img_array[22+cnt1][10+cnt2];\
					producted_1[67] <= in_img_array[22+cnt1][11+cnt2];\
					producted_1[68] <= in_img_array[22+cnt1][12+cnt2];\
					producted_1[69] <= in_img_array[22+cnt1][13+cnt2];\
					producted_1[70] <= in_img_array[22+cnt1][14+cnt2];\
					producted_1[71] <= in_img_array[22+cnt1][15+cnt2];\
					producted_1[72] <= in_img_array[22+cnt1][16+cnt2];\
					producted_1[73] <= in_img_array[22+cnt1][17+cnt2];\
					producted_1[74] <= in_img_array[22+cnt1][18+cnt2];\
					producted_1[75] <= in_img_array[22+cnt1][19+cnt2];\
					producted_1[76] <= in_img_array[22+cnt1][20+cnt2];\
					producted_1[77] <= in_img_array[22+cnt1][21+cnt2];\
					producted_1[78] <= in_img_array[22+cnt1][22+cnt2];\
					producted_1[79] <= in_img_array[22+cnt1][23+cnt2];\
					producted_1[80] <= in_img_array[22+cnt1][24+cnt2];\
					producted_1[81] <= in_img_array[22+cnt1][25+cnt2];\
					producted_1[82] <= in_img_array[22+cnt1][26+cnt2];\
					producted_1[83] <= in_img_array[22+cnt1][27+cnt2];\
					producted_1[84] <= in_img_array[23+cnt1][0+cnt2];\
					producted_1[85] <= in_img_array[23+cnt1][1+cnt2];\
					producted_1[86] <= in_img_array[23+cnt1][2+cnt2];\
					producted_1[87] <= in_img_array[23+cnt1][3+cnt2];\
					producted_1[88] <= in_img_array[23+cnt1][4+cnt2];\
					producted_1[89] <= in_img_array[23+cnt1][5+cnt2];\
					producted_1[90] <= in_img_array[23+cnt1][6+cnt2];\
					producted_1[91] <= in_img_array[23+cnt1][7+cnt2];\
					producted_1[92] <= in_img_array[23+cnt1][8+cnt2];\
					producted_1[93] <= in_img_array[23+cnt1][9+cnt2];\
					producted_1[94] <= in_img_array[23+cnt1][10+cnt2];\
					producted_1[95] <= in_img_array[23+cnt1][11+cnt2];\
					producted_1[96] <= in_img_array[23+cnt1][12+cnt2];\
					producted_1[97] <= in_img_array[23+cnt1][13+cnt2];\
					producted_1[98] <= in_img_array[23+cnt1][14+cnt2];\
					producted_1[99] <= in_img_array[23+cnt1][15+cnt2];\
					producted_1[100] <= in_img_array[23+cnt1][16+cnt2];\
					producted_1[101] <= in_img_array[23+cnt1][17+cnt2];\
					producted_1[102] <= in_img_array[23+cnt1][18+cnt2];\
					producted_1[103] <= in_img_array[23+cnt1][19+cnt2];\
					producted_1[104] <= in_img_array[23+cnt1][20+cnt2];\
					producted_1[105] <= in_img_array[23+cnt1][21+cnt2];\
					producted_1[106] <= in_img_array[23+cnt1][22+cnt2];\
					producted_1[107] <= in_img_array[23+cnt1][23+cnt2];\
					producted_1[108] <= in_img_array[23+cnt1][24+cnt2];\
					producted_1[109] <= in_img_array[23+cnt1][25+cnt2];\
					producted_1[110] <= in_img_array[23+cnt1][26+cnt2];\
					producted_1[111] <= in_img_array[23+cnt1][27+cnt2];\
                end\
            end\
            CONV1_1_7,CONV1_2_7,CONV1_3_7,CONV1_4_7,CONV1_5_7,CONV1_6_7:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_1[0] <= in_img_array[24+cnt1][0+cnt2];\
					producted_1[1] <= in_img_array[24+cnt1][1+cnt2];\
					producted_1[2] <= in_img_array[24+cnt1][2+cnt2];\
					producted_1[3] <= in_img_array[24+cnt1][3+cnt2];\
					producted_1[4] <= in_img_array[24+cnt1][4+cnt2];\
					producted_1[5] <= in_img_array[24+cnt1][5+cnt2];\
					producted_1[6] <= in_img_array[24+cnt1][6+cnt2];\
					producted_1[7] <= in_img_array[24+cnt1][7+cnt2];\
					producted_1[8] <= in_img_array[24+cnt1][8+cnt2];\
					producted_1[9] <= in_img_array[24+cnt1][9+cnt2];\
					producted_1[10] <= in_img_array[24+cnt1][10+cnt2];\
					producted_1[11] <= in_img_array[24+cnt1][11+cnt2];\
					producted_1[12] <= in_img_array[24+cnt1][12+cnt2];\
					producted_1[13] <= in_img_array[24+cnt1][13+cnt2];\
					producted_1[14] <= in_img_array[24+cnt1][14+cnt2];\
					producted_1[15] <= in_img_array[24+cnt1][15+cnt2];\
					producted_1[16] <= in_img_array[24+cnt1][16+cnt2];\
					producted_1[17] <= in_img_array[24+cnt1][17+cnt2];\
					producted_1[18] <= in_img_array[24+cnt1][18+cnt2];\
					producted_1[19] <= in_img_array[24+cnt1][19+cnt2];\
					producted_1[20] <= in_img_array[24+cnt1][20+cnt2];\
					producted_1[21] <= in_img_array[24+cnt1][21+cnt2];\
					producted_1[22] <= in_img_array[24+cnt1][22+cnt2];\
					producted_1[23] <= in_img_array[24+cnt1][23+cnt2];\
					producted_1[24] <= in_img_array[24+cnt1][24+cnt2];\
					producted_1[25] <= in_img_array[24+cnt1][25+cnt2];\
					producted_1[26] <= in_img_array[24+cnt1][26+cnt2];\
					producted_1[27] <= in_img_array[24+cnt1][27+cnt2];\
					producted_1[28] <= in_img_array[25+cnt1][0+cnt2];\
					producted_1[29] <= in_img_array[25+cnt1][1+cnt2];\
					producted_1[30] <= in_img_array[25+cnt1][2+cnt2];\
					producted_1[31] <= in_img_array[25+cnt1][3+cnt2];\
					producted_1[32] <= in_img_array[25+cnt1][4+cnt2];\
					producted_1[33] <= in_img_array[25+cnt1][5+cnt2];\
					producted_1[34] <= in_img_array[25+cnt1][6+cnt2];\
					producted_1[35] <= in_img_array[25+cnt1][7+cnt2];\
					producted_1[36] <= in_img_array[25+cnt1][8+cnt2];\
					producted_1[37] <= in_img_array[25+cnt1][9+cnt2];\
					producted_1[38] <= in_img_array[25+cnt1][10+cnt2];\
					producted_1[39] <= in_img_array[25+cnt1][11+cnt2];\
					producted_1[40] <= in_img_array[25+cnt1][12+cnt2];\
					producted_1[41] <= in_img_array[25+cnt1][13+cnt2];\
					producted_1[42] <= in_img_array[25+cnt1][14+cnt2];\
					producted_1[43] <= in_img_array[25+cnt1][15+cnt2];\
					producted_1[44] <= in_img_array[25+cnt1][16+cnt2];\
					producted_1[45] <= in_img_array[25+cnt1][17+cnt2];\
					producted_1[46] <= in_img_array[25+cnt1][18+cnt2];\
					producted_1[47] <= in_img_array[25+cnt1][19+cnt2];\
					producted_1[48] <= in_img_array[25+cnt1][20+cnt2];\
					producted_1[49] <= in_img_array[25+cnt1][21+cnt2];\
					producted_1[50] <= in_img_array[25+cnt1][22+cnt2];\
					producted_1[51] <= in_img_array[25+cnt1][23+cnt2];\
					producted_1[52] <= in_img_array[25+cnt1][24+cnt2];\
					producted_1[53] <= in_img_array[25+cnt1][25+cnt2];\
					producted_1[54] <= in_img_array[25+cnt1][26+cnt2];\
					producted_1[55] <= in_img_array[25+cnt1][27+cnt2];\
					producted_1[56] <= in_img_array[26+cnt1][0+cnt2];\
					producted_1[57] <= in_img_array[26+cnt1][1+cnt2];\
					producted_1[58] <= in_img_array[26+cnt1][2+cnt2];\
					producted_1[59] <= in_img_array[26+cnt1][3+cnt2];\
					producted_1[60] <= in_img_array[26+cnt1][4+cnt2];\
					producted_1[61] <= in_img_array[26+cnt1][5+cnt2];\
					producted_1[62] <= in_img_array[26+cnt1][6+cnt2];\
					producted_1[63] <= in_img_array[26+cnt1][7+cnt2];\
					producted_1[64] <= in_img_array[26+cnt1][8+cnt2];\
					producted_1[65] <= in_img_array[26+cnt1][9+cnt2];\
					producted_1[66] <= in_img_array[26+cnt1][10+cnt2];\
					producted_1[67] <= in_img_array[26+cnt1][11+cnt2];\
					producted_1[68] <= in_img_array[26+cnt1][12+cnt2];\
					producted_1[69] <= in_img_array[26+cnt1][13+cnt2];\
					producted_1[70] <= in_img_array[26+cnt1][14+cnt2];\
					producted_1[71] <= in_img_array[26+cnt1][15+cnt2];\
					producted_1[72] <= in_img_array[26+cnt1][16+cnt2];\
					producted_1[73] <= in_img_array[26+cnt1][17+cnt2];\
					producted_1[74] <= in_img_array[26+cnt1][18+cnt2];\
					producted_1[75] <= in_img_array[26+cnt1][19+cnt2];\
					producted_1[76] <= in_img_array[26+cnt1][20+cnt2];\
					producted_1[77] <= in_img_array[26+cnt1][21+cnt2];\
					producted_1[78] <= in_img_array[26+cnt1][22+cnt2];\
					producted_1[79] <= in_img_array[26+cnt1][23+cnt2];\
					producted_1[80] <= in_img_array[26+cnt1][24+cnt2];\
					producted_1[81] <= in_img_array[26+cnt1][25+cnt2];\
					producted_1[82] <= in_img_array[26+cnt1][26+cnt2];\
					producted_1[83] <= in_img_array[26+cnt1][27+cnt2];\
					producted_1[84] <= in_img_array[27+cnt1][0+cnt2];\
					producted_1[85] <= in_img_array[27+cnt1][1+cnt2];\
					producted_1[86] <= in_img_array[27+cnt1][2+cnt2];\
					producted_1[87] <= in_img_array[27+cnt1][3+cnt2];\
					producted_1[88] <= in_img_array[27+cnt1][4+cnt2];\
					producted_1[89] <= in_img_array[27+cnt1][5+cnt2];\
					producted_1[90] <= in_img_array[27+cnt1][6+cnt2];\
					producted_1[91] <= in_img_array[27+cnt1][7+cnt2];\
					producted_1[92] <= in_img_array[27+cnt1][8+cnt2];\
					producted_1[93] <= in_img_array[27+cnt1][9+cnt2];\
					producted_1[94] <= in_img_array[27+cnt1][10+cnt2];\
					producted_1[95] <= in_img_array[27+cnt1][11+cnt2];\
					producted_1[96] <= in_img_array[27+cnt1][12+cnt2];\
					producted_1[97] <= in_img_array[27+cnt1][13+cnt2];\
					producted_1[98] <= in_img_array[27+cnt1][14+cnt2];\
					producted_1[99] <= in_img_array[27+cnt1][15+cnt2];\
					producted_1[100] <= in_img_array[27+cnt1][16+cnt2];\
					producted_1[101] <= in_img_array[27+cnt1][17+cnt2];\
					producted_1[102] <= in_img_array[27+cnt1][18+cnt2];\
					producted_1[103] <= in_img_array[27+cnt1][19+cnt2];\
					producted_1[104] <= in_img_array[27+cnt1][20+cnt2];\
					producted_1[105] <= in_img_array[27+cnt1][21+cnt2];\
					producted_1[106] <= in_img_array[27+cnt1][22+cnt2];\
					producted_1[107] <= in_img_array[27+cnt1][23+cnt2];\
					producted_1[108] <= in_img_array[27+cnt1][24+cnt2];\
					producted_1[109] <= in_img_array[27+cnt1][25+cnt2];\
					producted_1[110] <= in_img_array[27+cnt1][26+cnt2];\
					producted_1[111] <= in_img_array[27+cnt1][27+cnt2];\
                end\
            end\
            CONV2_1_1,CONV2_2_1,CONV2_3_1,CONV2_4_1,CONV2_5_1,CONV2_6_1:begin\
				producted_1[0] <= conv1_result[0][0+cnt1][0+cnt2];\
				producted_1[1] <= conv1_result[0][0+cnt1][1+cnt2];\
				producted_1[2] <= conv1_result[0][0+cnt1][2+cnt2];\
				producted_1[3] <= conv1_result[0][0+cnt1][3+cnt2];\
				producted_1[4] <= conv1_result[0][0+cnt1][4+cnt2];\
				producted_1[5] <= conv1_result[0][0+cnt1][5+cnt2];\
				producted_1[6] <= conv1_result[0][0+cnt1][6+cnt2];\
				producted_1[7] <= conv1_result[0][0+cnt1][7+cnt2];\
				producted_1[8] <= conv1_result[0][0+cnt1][8+cnt2];\
				producted_1[9] <= conv1_result[0][0+cnt1][9+cnt2];\
				producted_1[10] <= conv1_result[0][1+cnt1][0+cnt2];\
				producted_1[11] <= conv1_result[0][1+cnt1][1+cnt2];\
				producted_1[12] <= conv1_result[0][1+cnt1][2+cnt2];\
				producted_1[13] <= conv1_result[0][1+cnt1][3+cnt2];\
				producted_1[14] <= conv1_result[0][1+cnt1][4+cnt2];\
				producted_1[15] <= conv1_result[0][1+cnt1][5+cnt2];\
				producted_1[16] <= conv1_result[0][1+cnt1][6+cnt2];\
				producted_1[17] <= conv1_result[0][1+cnt1][7+cnt2];\
				producted_1[18] <= conv1_result[0][1+cnt1][8+cnt2];\
				producted_1[19] <= conv1_result[0][1+cnt1][9+cnt2];\
				producted_1[20] <= conv1_result[0][2+cnt1][0+cnt2];\
				producted_1[21] <= conv1_result[0][2+cnt1][1+cnt2];\
				producted_1[22] <= conv1_result[0][2+cnt1][2+cnt2];\
				producted_1[23] <= conv1_result[0][2+cnt1][3+cnt2];\
				producted_1[24] <= conv1_result[0][2+cnt1][4+cnt2];\
				producted_1[25] <= conv1_result[0][2+cnt1][5+cnt2];\
				producted_1[26] <= conv1_result[0][2+cnt1][6+cnt2];\
				producted_1[27] <= conv1_result[0][2+cnt1][7+cnt2];\
				producted_1[28] <= conv1_result[0][2+cnt1][8+cnt2];\
				producted_1[29] <= conv1_result[0][2+cnt1][9+cnt2];\
				producted_1[30] <= conv1_result[0][3+cnt1][0+cnt2];\
				producted_1[31] <= conv1_result[0][3+cnt1][1+cnt2];\
				producted_1[32] <= conv1_result[0][3+cnt1][2+cnt2];\
				producted_1[33] <= conv1_result[0][3+cnt1][3+cnt2];\
				producted_1[34] <= conv1_result[0][3+cnt1][4+cnt2];\
				producted_1[35] <= conv1_result[0][3+cnt1][5+cnt2];\
				producted_1[36] <= conv1_result[0][3+cnt1][6+cnt2];\
				producted_1[37] <= conv1_result[0][3+cnt1][7+cnt2];\
				producted_1[38] <= conv1_result[0][3+cnt1][8+cnt2];\
				producted_1[39] <= conv1_result[0][3+cnt1][9+cnt2];\
				producted_1[40] <= conv1_result[0][4+cnt1][0+cnt2];\
				producted_1[41] <= conv1_result[0][4+cnt1][1+cnt2];\
				producted_1[42] <= conv1_result[0][4+cnt1][2+cnt2];\
				producted_1[43] <= conv1_result[0][4+cnt1][3+cnt2];\
				producted_1[44] <= conv1_result[0][4+cnt1][4+cnt2];\
				producted_1[45] <= conv1_result[0][4+cnt1][5+cnt2];\
				producted_1[46] <= conv1_result[0][4+cnt1][6+cnt2];\
				producted_1[47] <= conv1_result[0][4+cnt1][7+cnt2];\
				producted_1[48] <= conv1_result[0][4+cnt1][8+cnt2];\
				producted_1[49] <= conv1_result[0][4+cnt1][9+cnt2];\
				producted_1[50] <= conv1_result[0][5+cnt1][0+cnt2];\
				producted_1[51] <= conv1_result[0][5+cnt1][1+cnt2];\
				producted_1[52] <= conv1_result[0][5+cnt1][2+cnt2];\
				producted_1[53] <= conv1_result[0][5+cnt1][3+cnt2];\
				producted_1[54] <= conv1_result[0][5+cnt1][4+cnt2];\
				producted_1[55] <= conv1_result[0][5+cnt1][5+cnt2];\
				producted_1[56] <= conv1_result[0][5+cnt1][6+cnt2];\
				producted_1[57] <= conv1_result[0][5+cnt1][7+cnt2];\
				producted_1[58] <= conv1_result[0][5+cnt1][8+cnt2];\
				producted_1[59] <= conv1_result[0][5+cnt1][9+cnt2];\
				producted_1[60] <= conv1_result[0][6+cnt1][0+cnt2];\
				producted_1[61] <= conv1_result[0][6+cnt1][1+cnt2];\
				producted_1[62] <= conv1_result[0][6+cnt1][2+cnt2];\
				producted_1[63] <= conv1_result[0][6+cnt1][3+cnt2];\
				producted_1[64] <= conv1_result[0][6+cnt1][4+cnt2];\
				producted_1[65] <= conv1_result[0][6+cnt1][5+cnt2];\
				producted_1[66] <= conv1_result[0][6+cnt1][6+cnt2];\
				producted_1[67] <= conv1_result[0][6+cnt1][7+cnt2];\
				producted_1[68] <= conv1_result[0][6+cnt1][8+cnt2];\
				producted_1[69] <= conv1_result[0][6+cnt1][9+cnt2];\
				producted_1[70] <= conv1_result[0][7+cnt1][0+cnt2];\
				producted_1[71] <= conv1_result[0][7+cnt1][1+cnt2];\
				producted_1[72] <= conv1_result[0][7+cnt1][2+cnt2];\
				producted_1[73] <= conv1_result[0][7+cnt1][3+cnt2];\
				producted_1[74] <= conv1_result[0][7+cnt1][4+cnt2];\
				producted_1[75] <= conv1_result[0][7+cnt1][5+cnt2];\
				producted_1[76] <= conv1_result[0][7+cnt1][6+cnt2];\
				producted_1[77] <= conv1_result[0][7+cnt1][7+cnt2];\
				producted_1[78] <= conv1_result[0][7+cnt1][8+cnt2];\
				producted_1[79] <= conv1_result[0][7+cnt1][9+cnt2];\
				producted_1[80] <= conv1_result[0][8+cnt1][0+cnt2];\
				producted_1[81] <= conv1_result[0][8+cnt1][1+cnt2];\
				producted_1[82] <= conv1_result[0][8+cnt1][2+cnt2];\
				producted_1[83] <= conv1_result[0][8+cnt1][3+cnt2];\
				producted_1[84] <= conv1_result[0][8+cnt1][4+cnt2];\
				producted_1[85] <= conv1_result[0][8+cnt1][5+cnt2];\
				producted_1[86] <= conv1_result[0][8+cnt1][6+cnt2];\
				producted_1[87] <= conv1_result[0][8+cnt1][7+cnt2];\
				producted_1[88] <= conv1_result[0][8+cnt1][8+cnt2];\
				producted_1[89] <= conv1_result[0][8+cnt1][9+cnt2];\
				producted_1[90] <= conv1_result[0][9+cnt1][0+cnt2];\
				producted_1[91] <= conv1_result[0][9+cnt1][1+cnt2];\
				producted_1[92] <= conv1_result[0][9+cnt1][2+cnt2];\
				producted_1[93] <= conv1_result[0][9+cnt1][3+cnt2];\
				producted_1[94] <= conv1_result[0][9+cnt1][4+cnt2];\
				producted_1[95] <= conv1_result[0][9+cnt1][5+cnt2];\
				producted_1[96] <= conv1_result[0][9+cnt1][6+cnt2];\
				producted_1[97] <= conv1_result[0][9+cnt1][7+cnt2];\
				producted_1[98] <= conv1_result[0][9+cnt1][8+cnt2];\
				producted_1[99] <= conv1_result[0][9+cnt1][9+cnt2];\
				producted_1[100] <= 18'd0;\
				producted_1[101] <= 18'd0;\
				producted_1[102] <= 18'd0;\
				producted_1[103] <= 18'd0;\
				producted_1[104] <= 18'd0;\
				producted_1[105] <= 18'd0;\
				producted_1[106] <= 18'd0;\
				producted_1[107] <= 18'd0;\
				producted_1[108] <= 18'd0;\
				producted_1[109] <= 18'd0;\
				producted_1[110] <= 18'd0;\
				producted_1[111] <= 18'd0;\
            end\
            CONV2_1_2,CONV2_2_2,CONV2_3_2,CONV2_4_2,CONV2_5_2,CONV2_6_2:begin\
				producted_1[0] <= conv1_result[1][0+cnt1][0+cnt2];\
				producted_1[1] <= conv1_result[1][0+cnt1][1+cnt2];\
				producted_1[2] <= conv1_result[1][0+cnt1][2+cnt2];\
				producted_1[3] <= conv1_result[1][0+cnt1][3+cnt2];\
				producted_1[4] <= conv1_result[1][0+cnt1][4+cnt2];\
				producted_1[5] <= conv1_result[1][0+cnt1][5+cnt2];\
				producted_1[6] <= conv1_result[1][0+cnt1][6+cnt2];\
				producted_1[7] <= conv1_result[1][0+cnt1][7+cnt2];\
				producted_1[8] <= conv1_result[1][0+cnt1][8+cnt2];\
				producted_1[9] <= conv1_result[1][0+cnt1][9+cnt2];\
				producted_1[10] <= conv1_result[1][1+cnt1][0+cnt2];\
				producted_1[11] <= conv1_result[1][1+cnt1][1+cnt2];\
				producted_1[12] <= conv1_result[1][1+cnt1][2+cnt2];\
				producted_1[13] <= conv1_result[1][1+cnt1][3+cnt2];\
				producted_1[14] <= conv1_result[1][1+cnt1][4+cnt2];\
				producted_1[15] <= conv1_result[1][1+cnt1][5+cnt2];\
				producted_1[16] <= conv1_result[1][1+cnt1][6+cnt2];\
				producted_1[17] <= conv1_result[1][1+cnt1][7+cnt2];\
				producted_1[18] <= conv1_result[1][1+cnt1][8+cnt2];\
				producted_1[19] <= conv1_result[1][1+cnt1][9+cnt2];\
				producted_1[20] <= conv1_result[1][2+cnt1][0+cnt2];\
				producted_1[21] <= conv1_result[1][2+cnt1][1+cnt2];\
				producted_1[22] <= conv1_result[1][2+cnt1][2+cnt2];\
				producted_1[23] <= conv1_result[1][2+cnt1][3+cnt2];\
				producted_1[24] <= conv1_result[1][2+cnt1][4+cnt2];\
				producted_1[25] <= conv1_result[1][2+cnt1][5+cnt2];\
				producted_1[26] <= conv1_result[1][2+cnt1][6+cnt2];\
				producted_1[27] <= conv1_result[1][2+cnt1][7+cnt2];\
				producted_1[28] <= conv1_result[1][2+cnt1][8+cnt2];\
				producted_1[29] <= conv1_result[1][2+cnt1][9+cnt2];\
				producted_1[30] <= conv1_result[1][3+cnt1][0+cnt2];\
				producted_1[31] <= conv1_result[1][3+cnt1][1+cnt2];\
				producted_1[32] <= conv1_result[1][3+cnt1][2+cnt2];\
				producted_1[33] <= conv1_result[1][3+cnt1][3+cnt2];\
				producted_1[34] <= conv1_result[1][3+cnt1][4+cnt2];\
				producted_1[35] <= conv1_result[1][3+cnt1][5+cnt2];\
				producted_1[36] <= conv1_result[1][3+cnt1][6+cnt2];\
				producted_1[37] <= conv1_result[1][3+cnt1][7+cnt2];\
				producted_1[38] <= conv1_result[1][3+cnt1][8+cnt2];\
				producted_1[39] <= conv1_result[1][3+cnt1][9+cnt2];\
				producted_1[40] <= conv1_result[1][4+cnt1][0+cnt2];\
				producted_1[41] <= conv1_result[1][4+cnt1][1+cnt2];\
				producted_1[42] <= conv1_result[1][4+cnt1][2+cnt2];\
				producted_1[43] <= conv1_result[1][4+cnt1][3+cnt2];\
				producted_1[44] <= conv1_result[1][4+cnt1][4+cnt2];\
				producted_1[45] <= conv1_result[1][4+cnt1][5+cnt2];\
				producted_1[46] <= conv1_result[1][4+cnt1][6+cnt2];\
				producted_1[47] <= conv1_result[1][4+cnt1][7+cnt2];\
				producted_1[48] <= conv1_result[1][4+cnt1][8+cnt2];\
				producted_1[49] <= conv1_result[1][4+cnt1][9+cnt2];\
				producted_1[50] <= conv1_result[1][5+cnt1][0+cnt2];\
				producted_1[51] <= conv1_result[1][5+cnt1][1+cnt2];\
				producted_1[52] <= conv1_result[1][5+cnt1][2+cnt2];\
				producted_1[53] <= conv1_result[1][5+cnt1][3+cnt2];\
				producted_1[54] <= conv1_result[1][5+cnt1][4+cnt2];\
				producted_1[55] <= conv1_result[1][5+cnt1][5+cnt2];\
				producted_1[56] <= conv1_result[1][5+cnt1][6+cnt2];\
				producted_1[57] <= conv1_result[1][5+cnt1][7+cnt2];\
				producted_1[58] <= conv1_result[1][5+cnt1][8+cnt2];\
				producted_1[59] <= conv1_result[1][5+cnt1][9+cnt2];\
				producted_1[60] <= conv1_result[1][6+cnt1][0+cnt2];\
				producted_1[61] <= conv1_result[1][6+cnt1][1+cnt2];\
				producted_1[62] <= conv1_result[1][6+cnt1][2+cnt2];\
				producted_1[63] <= conv1_result[1][6+cnt1][3+cnt2];\
				producted_1[64] <= conv1_result[1][6+cnt1][4+cnt2];\
				producted_1[65] <= conv1_result[1][6+cnt1][5+cnt2];\
				producted_1[66] <= conv1_result[1][6+cnt1][6+cnt2];\
				producted_1[67] <= conv1_result[1][6+cnt1][7+cnt2];\
				producted_1[68] <= conv1_result[1][6+cnt1][8+cnt2];\
				producted_1[69] <= conv1_result[1][6+cnt1][9+cnt2];\
				producted_1[70] <= conv1_result[1][7+cnt1][0+cnt2];\
				producted_1[71] <= conv1_result[1][7+cnt1][1+cnt2];\
				producted_1[72] <= conv1_result[1][7+cnt1][2+cnt2];\
				producted_1[73] <= conv1_result[1][7+cnt1][3+cnt2];\
				producted_1[74] <= conv1_result[1][7+cnt1][4+cnt2];\
				producted_1[75] <= conv1_result[1][7+cnt1][5+cnt2];\
				producted_1[76] <= conv1_result[1][7+cnt1][6+cnt2];\
				producted_1[77] <= conv1_result[1][7+cnt1][7+cnt2];\
				producted_1[78] <= conv1_result[1][7+cnt1][8+cnt2];\
				producted_1[79] <= conv1_result[1][7+cnt1][9+cnt2];\
				producted_1[80] <= conv1_result[1][8+cnt1][0+cnt2];\
				producted_1[81] <= conv1_result[1][8+cnt1][1+cnt2];\
				producted_1[82] <= conv1_result[1][8+cnt1][2+cnt2];\
				producted_1[83] <= conv1_result[1][8+cnt1][3+cnt2];\
				producted_1[84] <= conv1_result[1][8+cnt1][4+cnt2];\
				producted_1[85] <= conv1_result[1][8+cnt1][5+cnt2];\
				producted_1[86] <= conv1_result[1][8+cnt1][6+cnt2];\
				producted_1[87] <= conv1_result[1][8+cnt1][7+cnt2];\
				producted_1[88] <= conv1_result[1][8+cnt1][8+cnt2];\
				producted_1[89] <= conv1_result[1][8+cnt1][9+cnt2];\
				producted_1[90] <= conv1_result[1][9+cnt1][0+cnt2];\
				producted_1[91] <= conv1_result[1][9+cnt1][1+cnt2];\
				producted_1[92] <= conv1_result[1][9+cnt1][2+cnt2];\
				producted_1[93] <= conv1_result[1][9+cnt1][3+cnt2];\
				producted_1[94] <= conv1_result[1][9+cnt1][4+cnt2];\
				producted_1[95] <= conv1_result[1][9+cnt1][5+cnt2];\
				producted_1[96] <= conv1_result[1][9+cnt1][6+cnt2];\
				producted_1[97] <= conv1_result[1][9+cnt1][7+cnt2];\
				producted_1[98] <= conv1_result[1][9+cnt1][8+cnt2];\
				producted_1[99] <= conv1_result[1][9+cnt1][9+cnt2];\
				producted_1[100] <= 18'd0;\
				producted_1[101] <= 18'd0;\
				producted_1[102] <= 18'd0;\
				producted_1[103] <= 18'd0;\
				producted_1[104] <= 18'd0;\
				producted_1[105] <= 18'd0;\
				producted_1[106] <= 18'd0;\
				producted_1[107] <= 18'd0;\
				producted_1[108] <= 18'd0;\
				producted_1[109] <= 18'd0;\
				producted_1[110] <= 18'd0;\
				producted_1[111] <= 18'd0;\
            end\
            CONV2_1_3,CONV2_2_3,CONV2_3_3,CONV2_4_3,CONV2_5_3,CONV2_6_3:begin\
				producted_1[0] <= conv1_result[2][0+cnt1][0+cnt2];\
				producted_1[1] <= conv1_result[2][0+cnt1][1+cnt2];\
				producted_1[2] <= conv1_result[2][0+cnt1][2+cnt2];\
				producted_1[3] <= conv1_result[2][0+cnt1][3+cnt2];\
				producted_1[4] <= conv1_result[2][0+cnt1][4+cnt2];\
				producted_1[5] <= conv1_result[2][0+cnt1][5+cnt2];\
				producted_1[6] <= conv1_result[2][0+cnt1][6+cnt2];\
				producted_1[7] <= conv1_result[2][0+cnt1][7+cnt2];\
				producted_1[8] <= conv1_result[2][0+cnt1][8+cnt2];\
				producted_1[9] <= conv1_result[2][0+cnt1][9+cnt2];\
				producted_1[10] <= conv1_result[2][1+cnt1][0+cnt2];\
				producted_1[11] <= conv1_result[2][1+cnt1][1+cnt2];\
				producted_1[12] <= conv1_result[2][1+cnt1][2+cnt2];\
				producted_1[13] <= conv1_result[2][1+cnt1][3+cnt2];\
				producted_1[14] <= conv1_result[2][1+cnt1][4+cnt2];\
				producted_1[15] <= conv1_result[2][1+cnt1][5+cnt2];\
				producted_1[16] <= conv1_result[2][1+cnt1][6+cnt2];\
				producted_1[17] <= conv1_result[2][1+cnt1][7+cnt2];\
				producted_1[18] <= conv1_result[2][1+cnt1][8+cnt2];\
				producted_1[19] <= conv1_result[2][1+cnt1][9+cnt2];\
				producted_1[20] <= conv1_result[2][2+cnt1][0+cnt2];\
				producted_1[21] <= conv1_result[2][2+cnt1][1+cnt2];\
				producted_1[22] <= conv1_result[2][2+cnt1][2+cnt2];\
				producted_1[23] <= conv1_result[2][2+cnt1][3+cnt2];\
				producted_1[24] <= conv1_result[2][2+cnt1][4+cnt2];\
				producted_1[25] <= conv1_result[2][2+cnt1][5+cnt2];\
				producted_1[26] <= conv1_result[2][2+cnt1][6+cnt2];\
				producted_1[27] <= conv1_result[2][2+cnt1][7+cnt2];\
				producted_1[28] <= conv1_result[2][2+cnt1][8+cnt2];\
				producted_1[29] <= conv1_result[2][2+cnt1][9+cnt2];\
				producted_1[30] <= conv1_result[2][3+cnt1][0+cnt2];\
				producted_1[31] <= conv1_result[2][3+cnt1][1+cnt2];\
				producted_1[32] <= conv1_result[2][3+cnt1][2+cnt2];\
				producted_1[33] <= conv1_result[2][3+cnt1][3+cnt2];\
				producted_1[34] <= conv1_result[2][3+cnt1][4+cnt2];\
				producted_1[35] <= conv1_result[2][3+cnt1][5+cnt2];\
				producted_1[36] <= conv1_result[2][3+cnt1][6+cnt2];\
				producted_1[37] <= conv1_result[2][3+cnt1][7+cnt2];\
				producted_1[38] <= conv1_result[2][3+cnt1][8+cnt2];\
				producted_1[39] <= conv1_result[2][3+cnt1][9+cnt2];\
				producted_1[40] <= conv1_result[2][4+cnt1][0+cnt2];\
				producted_1[41] <= conv1_result[2][4+cnt1][1+cnt2];\
				producted_1[42] <= conv1_result[2][4+cnt1][2+cnt2];\
				producted_1[43] <= conv1_result[2][4+cnt1][3+cnt2];\
				producted_1[44] <= conv1_result[2][4+cnt1][4+cnt2];\
				producted_1[45] <= conv1_result[2][4+cnt1][5+cnt2];\
				producted_1[46] <= conv1_result[2][4+cnt1][6+cnt2];\
				producted_1[47] <= conv1_result[2][4+cnt1][7+cnt2];\
				producted_1[48] <= conv1_result[2][4+cnt1][8+cnt2];\
				producted_1[49] <= conv1_result[2][4+cnt1][9+cnt2];\
				producted_1[50] <= conv1_result[2][5+cnt1][0+cnt2];\
				producted_1[51] <= conv1_result[2][5+cnt1][1+cnt2];\
				producted_1[52] <= conv1_result[2][5+cnt1][2+cnt2];\
				producted_1[53] <= conv1_result[2][5+cnt1][3+cnt2];\
				producted_1[54] <= conv1_result[2][5+cnt1][4+cnt2];\
				producted_1[55] <= conv1_result[2][5+cnt1][5+cnt2];\
				producted_1[56] <= conv1_result[2][5+cnt1][6+cnt2];\
				producted_1[57] <= conv1_result[2][5+cnt1][7+cnt2];\
				producted_1[58] <= conv1_result[2][5+cnt1][8+cnt2];\
				producted_1[59] <= conv1_result[2][5+cnt1][9+cnt2];\
				producted_1[60] <= conv1_result[2][6+cnt1][0+cnt2];\
				producted_1[61] <= conv1_result[2][6+cnt1][1+cnt2];\
				producted_1[62] <= conv1_result[2][6+cnt1][2+cnt2];\
				producted_1[63] <= conv1_result[2][6+cnt1][3+cnt2];\
				producted_1[64] <= conv1_result[2][6+cnt1][4+cnt2];\
				producted_1[65] <= conv1_result[2][6+cnt1][5+cnt2];\
				producted_1[66] <= conv1_result[2][6+cnt1][6+cnt2];\
				producted_1[67] <= conv1_result[2][6+cnt1][7+cnt2];\
				producted_1[68] <= conv1_result[2][6+cnt1][8+cnt2];\
				producted_1[69] <= conv1_result[2][6+cnt1][9+cnt2];\
				producted_1[70] <= conv1_result[2][7+cnt1][0+cnt2];\
				producted_1[71] <= conv1_result[2][7+cnt1][1+cnt2];\
				producted_1[72] <= conv1_result[2][7+cnt1][2+cnt2];\
				producted_1[73] <= conv1_result[2][7+cnt1][3+cnt2];\
				producted_1[74] <= conv1_result[2][7+cnt1][4+cnt2];\
				producted_1[75] <= conv1_result[2][7+cnt1][5+cnt2];\
				producted_1[76] <= conv1_result[2][7+cnt1][6+cnt2];\
				producted_1[77] <= conv1_result[2][7+cnt1][7+cnt2];\
				producted_1[78] <= conv1_result[2][7+cnt1][8+cnt2];\
				producted_1[79] <= conv1_result[2][7+cnt1][9+cnt2];\
				producted_1[80] <= conv1_result[2][8+cnt1][0+cnt2];\
				producted_1[81] <= conv1_result[2][8+cnt1][1+cnt2];\
				producted_1[82] <= conv1_result[2][8+cnt1][2+cnt2];\
				producted_1[83] <= conv1_result[2][8+cnt1][3+cnt2];\
				producted_1[84] <= conv1_result[2][8+cnt1][4+cnt2];\
				producted_1[85] <= conv1_result[2][8+cnt1][5+cnt2];\
				producted_1[86] <= conv1_result[2][8+cnt1][6+cnt2];\
				producted_1[87] <= conv1_result[2][8+cnt1][7+cnt2];\
				producted_1[88] <= conv1_result[2][8+cnt1][8+cnt2];\
				producted_1[89] <= conv1_result[2][8+cnt1][9+cnt2];\
				producted_1[90] <= conv1_result[2][9+cnt1][0+cnt2];\
				producted_1[91] <= conv1_result[2][9+cnt1][1+cnt2];\
				producted_1[92] <= conv1_result[2][9+cnt1][2+cnt2];\
				producted_1[93] <= conv1_result[2][9+cnt1][3+cnt2];\
				producted_1[94] <= conv1_result[2][9+cnt1][4+cnt2];\
				producted_1[95] <= conv1_result[2][9+cnt1][5+cnt2];\
				producted_1[96] <= conv1_result[2][9+cnt1][6+cnt2];\
				producted_1[97] <= conv1_result[2][9+cnt1][7+cnt2];\
				producted_1[98] <= conv1_result[2][9+cnt1][8+cnt2];\
				producted_1[99] <= conv1_result[2][9+cnt1][9+cnt2];\
				producted_1[100] <= 18'd0;\
				producted_1[101] <= 18'd0;\
				producted_1[102] <= 18'd0;\
				producted_1[103] <= 18'd0;\
				producted_1[104] <= 18'd0;\
				producted_1[105] <= 18'd0;\
				producted_1[106] <= 18'd0;\
				producted_1[107] <= 18'd0;\
				producted_1[108] <= 18'd0;\
				producted_1[109] <= 18'd0;\
				producted_1[110] <= 18'd0;\
				producted_1[111] <= 18'd0;\
            end\
            CONV2_1_4,CONV2_2_4,CONV2_3_4,CONV2_4_4,CONV2_5_4,CONV2_6_4:begin\
				producted_1[0] <= conv1_result[3][0+cnt1][0+cnt2];\
				producted_1[1] <= conv1_result[3][0+cnt1][1+cnt2];\
				producted_1[2] <= conv1_result[3][0+cnt1][2+cnt2];\
				producted_1[3] <= conv1_result[3][0+cnt1][3+cnt2];\
				producted_1[4] <= conv1_result[3][0+cnt1][4+cnt2];\
				producted_1[5] <= conv1_result[3][0+cnt1][5+cnt2];\
				producted_1[6] <= conv1_result[3][0+cnt1][6+cnt2];\
				producted_1[7] <= conv1_result[3][0+cnt1][7+cnt2];\
				producted_1[8] <= conv1_result[3][0+cnt1][8+cnt2];\
				producted_1[9] <= conv1_result[3][0+cnt1][9+cnt2];\
				producted_1[10] <= conv1_result[3][1+cnt1][0+cnt2];\
				producted_1[11] <= conv1_result[3][1+cnt1][1+cnt2];\
				producted_1[12] <= conv1_result[3][1+cnt1][2+cnt2];\
				producted_1[13] <= conv1_result[3][1+cnt1][3+cnt2];\
				producted_1[14] <= conv1_result[3][1+cnt1][4+cnt2];\
				producted_1[15] <= conv1_result[3][1+cnt1][5+cnt2];\
				producted_1[16] <= conv1_result[3][1+cnt1][6+cnt2];\
				producted_1[17] <= conv1_result[3][1+cnt1][7+cnt2];\
				producted_1[18] <= conv1_result[3][1+cnt1][8+cnt2];\
				producted_1[19] <= conv1_result[3][1+cnt1][9+cnt2];\
				producted_1[20] <= conv1_result[3][2+cnt1][0+cnt2];\
				producted_1[21] <= conv1_result[3][2+cnt1][1+cnt2];\
				producted_1[22] <= conv1_result[3][2+cnt1][2+cnt2];\
				producted_1[23] <= conv1_result[3][2+cnt1][3+cnt2];\
				producted_1[24] <= conv1_result[3][2+cnt1][4+cnt2];\
				producted_1[25] <= conv1_result[3][2+cnt1][5+cnt2];\
				producted_1[26] <= conv1_result[3][2+cnt1][6+cnt2];\
				producted_1[27] <= conv1_result[3][2+cnt1][7+cnt2];\
				producted_1[28] <= conv1_result[3][2+cnt1][8+cnt2];\
				producted_1[29] <= conv1_result[3][2+cnt1][9+cnt2];\
				producted_1[30] <= conv1_result[3][3+cnt1][0+cnt2];\
				producted_1[31] <= conv1_result[3][3+cnt1][1+cnt2];\
				producted_1[32] <= conv1_result[3][3+cnt1][2+cnt2];\
				producted_1[33] <= conv1_result[3][3+cnt1][3+cnt2];\
				producted_1[34] <= conv1_result[3][3+cnt1][4+cnt2];\
				producted_1[35] <= conv1_result[3][3+cnt1][5+cnt2];\
				producted_1[36] <= conv1_result[3][3+cnt1][6+cnt2];\
				producted_1[37] <= conv1_result[3][3+cnt1][7+cnt2];\
				producted_1[38] <= conv1_result[3][3+cnt1][8+cnt2];\
				producted_1[39] <= conv1_result[3][3+cnt1][9+cnt2];\
				producted_1[40] <= conv1_result[3][4+cnt1][0+cnt2];\
				producted_1[41] <= conv1_result[3][4+cnt1][1+cnt2];\
				producted_1[42] <= conv1_result[3][4+cnt1][2+cnt2];\
				producted_1[43] <= conv1_result[3][4+cnt1][3+cnt2];\
				producted_1[44] <= conv1_result[3][4+cnt1][4+cnt2];\
				producted_1[45] <= conv1_result[3][4+cnt1][5+cnt2];\
				producted_1[46] <= conv1_result[3][4+cnt1][6+cnt2];\
				producted_1[47] <= conv1_result[3][4+cnt1][7+cnt2];\
				producted_1[48] <= conv1_result[3][4+cnt1][8+cnt2];\
				producted_1[49] <= conv1_result[3][4+cnt1][9+cnt2];\
				producted_1[50] <= conv1_result[3][5+cnt1][0+cnt2];\
				producted_1[51] <= conv1_result[3][5+cnt1][1+cnt2];\
				producted_1[52] <= conv1_result[3][5+cnt1][2+cnt2];\
				producted_1[53] <= conv1_result[3][5+cnt1][3+cnt2];\
				producted_1[54] <= conv1_result[3][5+cnt1][4+cnt2];\
				producted_1[55] <= conv1_result[3][5+cnt1][5+cnt2];\
				producted_1[56] <= conv1_result[3][5+cnt1][6+cnt2];\
				producted_1[57] <= conv1_result[3][5+cnt1][7+cnt2];\
				producted_1[58] <= conv1_result[3][5+cnt1][8+cnt2];\
				producted_1[59] <= conv1_result[3][5+cnt1][9+cnt2];\
				producted_1[60] <= conv1_result[3][6+cnt1][0+cnt2];\
				producted_1[61] <= conv1_result[3][6+cnt1][1+cnt2];\
				producted_1[62] <= conv1_result[3][6+cnt1][2+cnt2];\
				producted_1[63] <= conv1_result[3][6+cnt1][3+cnt2];\
				producted_1[64] <= conv1_result[3][6+cnt1][4+cnt2];\
				producted_1[65] <= conv1_result[3][6+cnt1][5+cnt2];\
				producted_1[66] <= conv1_result[3][6+cnt1][6+cnt2];\
				producted_1[67] <= conv1_result[3][6+cnt1][7+cnt2];\
				producted_1[68] <= conv1_result[3][6+cnt1][8+cnt2];\
				producted_1[69] <= conv1_result[3][6+cnt1][9+cnt2];\
				producted_1[70] <= conv1_result[3][7+cnt1][0+cnt2];\
				producted_1[71] <= conv1_result[3][7+cnt1][1+cnt2];\
				producted_1[72] <= conv1_result[3][7+cnt1][2+cnt2];\
				producted_1[73] <= conv1_result[3][7+cnt1][3+cnt2];\
				producted_1[74] <= conv1_result[3][7+cnt1][4+cnt2];\
				producted_1[75] <= conv1_result[3][7+cnt1][5+cnt2];\
				producted_1[76] <= conv1_result[3][7+cnt1][6+cnt2];\
				producted_1[77] <= conv1_result[3][7+cnt1][7+cnt2];\
				producted_1[78] <= conv1_result[3][7+cnt1][8+cnt2];\
				producted_1[79] <= conv1_result[3][7+cnt1][9+cnt2];\
				producted_1[80] <= conv1_result[3][8+cnt1][0+cnt2];\
				producted_1[81] <= conv1_result[3][8+cnt1][1+cnt2];\
				producted_1[82] <= conv1_result[3][8+cnt1][2+cnt2];\
				producted_1[83] <= conv1_result[3][8+cnt1][3+cnt2];\
				producted_1[84] <= conv1_result[3][8+cnt1][4+cnt2];\
				producted_1[85] <= conv1_result[3][8+cnt1][5+cnt2];\
				producted_1[86] <= conv1_result[3][8+cnt1][6+cnt2];\
				producted_1[87] <= conv1_result[3][8+cnt1][7+cnt2];\
				producted_1[88] <= conv1_result[3][8+cnt1][8+cnt2];\
				producted_1[89] <= conv1_result[3][8+cnt1][9+cnt2];\
				producted_1[90] <= conv1_result[3][9+cnt1][0+cnt2];\
				producted_1[91] <= conv1_result[3][9+cnt1][1+cnt2];\
				producted_1[92] <= conv1_result[3][9+cnt1][2+cnt2];\
				producted_1[93] <= conv1_result[3][9+cnt1][3+cnt2];\
				producted_1[94] <= conv1_result[3][9+cnt1][4+cnt2];\
				producted_1[95] <= conv1_result[3][9+cnt1][5+cnt2];\
				producted_1[96] <= conv1_result[3][9+cnt1][6+cnt2];\
				producted_1[97] <= conv1_result[3][9+cnt1][7+cnt2];\
				producted_1[98] <= conv1_result[3][9+cnt1][8+cnt2];\
				producted_1[99] <= conv1_result[3][9+cnt1][9+cnt2];\
				producted_1[100] <= 18'd0;\
				producted_1[101] <= 18'd0;\
				producted_1[102] <= 18'd0;\
				producted_1[103] <= 18'd0;\
				producted_1[104] <= 18'd0;\
				producted_1[105] <= 18'd0;\
				producted_1[106] <= 18'd0;\
				producted_1[107] <= 18'd0;\
				producted_1[108] <= 18'd0;\
				producted_1[109] <= 18'd0;\
				producted_1[110] <= 18'd0;\
				producted_1[111] <= 18'd0;\
            end\
            CONV2_1_5,CONV2_2_5,CONV2_3_5,CONV2_4_5,CONV2_5_5,CONV2_6_5:begin\
				producted_1[0] <= conv1_result[4][0+cnt1][0+cnt2];\
				producted_1[1] <= conv1_result[4][0+cnt1][1+cnt2];\
				producted_1[2] <= conv1_result[4][0+cnt1][2+cnt2];\
				producted_1[3] <= conv1_result[4][0+cnt1][3+cnt2];\
				producted_1[4] <= conv1_result[4][0+cnt1][4+cnt2];\
				producted_1[5] <= conv1_result[4][0+cnt1][5+cnt2];\
				producted_1[6] <= conv1_result[4][0+cnt1][6+cnt2];\
				producted_1[7] <= conv1_result[4][0+cnt1][7+cnt2];\
				producted_1[8] <= conv1_result[4][0+cnt1][8+cnt2];\
				producted_1[9] <= conv1_result[4][0+cnt1][9+cnt2];\
				producted_1[10] <= conv1_result[4][1+cnt1][0+cnt2];\
				producted_1[11] <= conv1_result[4][1+cnt1][1+cnt2];\
				producted_1[12] <= conv1_result[4][1+cnt1][2+cnt2];\
				producted_1[13] <= conv1_result[4][1+cnt1][3+cnt2];\
				producted_1[14] <= conv1_result[4][1+cnt1][4+cnt2];\
				producted_1[15] <= conv1_result[4][1+cnt1][5+cnt2];\
				producted_1[16] <= conv1_result[4][1+cnt1][6+cnt2];\
				producted_1[17] <= conv1_result[4][1+cnt1][7+cnt2];\
				producted_1[18] <= conv1_result[4][1+cnt1][8+cnt2];\
				producted_1[19] <= conv1_result[4][1+cnt1][9+cnt2];\
				producted_1[20] <= conv1_result[4][2+cnt1][0+cnt2];\
				producted_1[21] <= conv1_result[4][2+cnt1][1+cnt2];\
				producted_1[22] <= conv1_result[4][2+cnt1][2+cnt2];\
				producted_1[23] <= conv1_result[4][2+cnt1][3+cnt2];\
				producted_1[24] <= conv1_result[4][2+cnt1][4+cnt2];\
				producted_1[25] <= conv1_result[4][2+cnt1][5+cnt2];\
				producted_1[26] <= conv1_result[4][2+cnt1][6+cnt2];\
				producted_1[27] <= conv1_result[4][2+cnt1][7+cnt2];\
				producted_1[28] <= conv1_result[4][2+cnt1][8+cnt2];\
				producted_1[29] <= conv1_result[4][2+cnt1][9+cnt2];\
				producted_1[30] <= conv1_result[4][3+cnt1][0+cnt2];\
				producted_1[31] <= conv1_result[4][3+cnt1][1+cnt2];\
				producted_1[32] <= conv1_result[4][3+cnt1][2+cnt2];\
				producted_1[33] <= conv1_result[4][3+cnt1][3+cnt2];\
				producted_1[34] <= conv1_result[4][3+cnt1][4+cnt2];\
				producted_1[35] <= conv1_result[4][3+cnt1][5+cnt2];\
				producted_1[36] <= conv1_result[4][3+cnt1][6+cnt2];\
				producted_1[37] <= conv1_result[4][3+cnt1][7+cnt2];\
				producted_1[38] <= conv1_result[4][3+cnt1][8+cnt2];\
				producted_1[39] <= conv1_result[4][3+cnt1][9+cnt2];\
				producted_1[40] <= conv1_result[4][4+cnt1][0+cnt2];\
				producted_1[41] <= conv1_result[4][4+cnt1][1+cnt2];\
				producted_1[42] <= conv1_result[4][4+cnt1][2+cnt2];\
				producted_1[43] <= conv1_result[4][4+cnt1][3+cnt2];\
				producted_1[44] <= conv1_result[4][4+cnt1][4+cnt2];\
				producted_1[45] <= conv1_result[4][4+cnt1][5+cnt2];\
				producted_1[46] <= conv1_result[4][4+cnt1][6+cnt2];\
				producted_1[47] <= conv1_result[4][4+cnt1][7+cnt2];\
				producted_1[48] <= conv1_result[4][4+cnt1][8+cnt2];\
				producted_1[49] <= conv1_result[4][4+cnt1][9+cnt2];\
				producted_1[50] <= conv1_result[4][5+cnt1][0+cnt2];\
				producted_1[51] <= conv1_result[4][5+cnt1][1+cnt2];\
				producted_1[52] <= conv1_result[4][5+cnt1][2+cnt2];\
				producted_1[53] <= conv1_result[4][5+cnt1][3+cnt2];\
				producted_1[54] <= conv1_result[4][5+cnt1][4+cnt2];\
				producted_1[55] <= conv1_result[4][5+cnt1][5+cnt2];\
				producted_1[56] <= conv1_result[4][5+cnt1][6+cnt2];\
				producted_1[57] <= conv1_result[4][5+cnt1][7+cnt2];\
				producted_1[58] <= conv1_result[4][5+cnt1][8+cnt2];\
				producted_1[59] <= conv1_result[4][5+cnt1][9+cnt2];\
				producted_1[60] <= conv1_result[4][6+cnt1][0+cnt2];\
				producted_1[61] <= conv1_result[4][6+cnt1][1+cnt2];\
				producted_1[62] <= conv1_result[4][6+cnt1][2+cnt2];\
				producted_1[63] <= conv1_result[4][6+cnt1][3+cnt2];\
				producted_1[64] <= conv1_result[4][6+cnt1][4+cnt2];\
				producted_1[65] <= conv1_result[4][6+cnt1][5+cnt2];\
				producted_1[66] <= conv1_result[4][6+cnt1][6+cnt2];\
				producted_1[67] <= conv1_result[4][6+cnt1][7+cnt2];\
				producted_1[68] <= conv1_result[4][6+cnt1][8+cnt2];\
				producted_1[69] <= conv1_result[4][6+cnt1][9+cnt2];\
				producted_1[70] <= conv1_result[4][7+cnt1][0+cnt2];\
				producted_1[71] <= conv1_result[4][7+cnt1][1+cnt2];\
				producted_1[72] <= conv1_result[4][7+cnt1][2+cnt2];\
				producted_1[73] <= conv1_result[4][7+cnt1][3+cnt2];\
				producted_1[74] <= conv1_result[4][7+cnt1][4+cnt2];\
				producted_1[75] <= conv1_result[4][7+cnt1][5+cnt2];\
				producted_1[76] <= conv1_result[4][7+cnt1][6+cnt2];\
				producted_1[77] <= conv1_result[4][7+cnt1][7+cnt2];\
				producted_1[78] <= conv1_result[4][7+cnt1][8+cnt2];\
				producted_1[79] <= conv1_result[4][7+cnt1][9+cnt2];\
				producted_1[80] <= conv1_result[4][8+cnt1][0+cnt2];\
				producted_1[81] <= conv1_result[4][8+cnt1][1+cnt2];\
				producted_1[82] <= conv1_result[4][8+cnt1][2+cnt2];\
				producted_1[83] <= conv1_result[4][8+cnt1][3+cnt2];\
				producted_1[84] <= conv1_result[4][8+cnt1][4+cnt2];\
				producted_1[85] <= conv1_result[4][8+cnt1][5+cnt2];\
				producted_1[86] <= conv1_result[4][8+cnt1][6+cnt2];\
				producted_1[87] <= conv1_result[4][8+cnt1][7+cnt2];\
				producted_1[88] <= conv1_result[4][8+cnt1][8+cnt2];\
				producted_1[89] <= conv1_result[4][8+cnt1][9+cnt2];\
				producted_1[90] <= conv1_result[4][9+cnt1][0+cnt2];\
				producted_1[91] <= conv1_result[4][9+cnt1][1+cnt2];\
				producted_1[92] <= conv1_result[4][9+cnt1][2+cnt2];\
				producted_1[93] <= conv1_result[4][9+cnt1][3+cnt2];\
				producted_1[94] <= conv1_result[4][9+cnt1][4+cnt2];\
				producted_1[95] <= conv1_result[4][9+cnt1][5+cnt2];\
				producted_1[96] <= conv1_result[4][9+cnt1][6+cnt2];\
				producted_1[97] <= conv1_result[4][9+cnt1][7+cnt2];\
				producted_1[98] <= conv1_result[4][9+cnt1][8+cnt2];\
				producted_1[99] <= conv1_result[4][9+cnt1][9+cnt2];\
				producted_1[100] <= 18'd0;\
				producted_1[101] <= 18'd0;\
				producted_1[102] <= 18'd0;\
				producted_1[103] <= 18'd0;\
				producted_1[104] <= 18'd0;\
				producted_1[105] <= 18'd0;\
				producted_1[106] <= 18'd0;\
				producted_1[107] <= 18'd0;\
				producted_1[108] <= 18'd0;\
				producted_1[109] <= 18'd0;\
				producted_1[110] <= 18'd0;\
				producted_1[111] <= 18'd0;\
            end\
            CONV2_1_6,CONV2_2_6,CONV2_3_6,CONV2_4_6,CONV2_5_6,CONV2_6_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_1[0] <= conv1_result[5][0+cnt1][0+cnt2];\
                    producted_1[1] <= conv1_result[5][0+cnt1][1+cnt2];\
                    producted_1[2] <= conv1_result[5][0+cnt1][2+cnt2];\
                    producted_1[3] <= conv1_result[5][0+cnt1][3+cnt2];\
                    producted_1[4] <= conv1_result[5][0+cnt1][4+cnt2];\
                    producted_1[5] <= conv1_result[5][0+cnt1][5+cnt2];\
                    producted_1[6] <= conv1_result[5][0+cnt1][6+cnt2];\
                    producted_1[7] <= conv1_result[5][0+cnt1][7+cnt2];\
                    producted_1[8] <= conv1_result[5][0+cnt1][8+cnt2];\
                    producted_1[9] <= conv1_result[5][0+cnt1][9+cnt2];\
                    producted_1[10] <= conv1_result[5][1+cnt1][0+cnt2];\
                    producted_1[11] <= conv1_result[5][1+cnt1][1+cnt2];\
                    producted_1[12] <= conv1_result[5][1+cnt1][2+cnt2];\
                    producted_1[13] <= conv1_result[5][1+cnt1][3+cnt2];\
                    producted_1[14] <= conv1_result[5][1+cnt1][4+cnt2];\
                    producted_1[15] <= conv1_result[5][1+cnt1][5+cnt2];\
                    producted_1[16] <= conv1_result[5][1+cnt1][6+cnt2];\
                    producted_1[17] <= conv1_result[5][1+cnt1][7+cnt2];\
                    producted_1[18] <= conv1_result[5][1+cnt1][8+cnt2];\
                    producted_1[19] <= conv1_result[5][1+cnt1][9+cnt2];\
                    producted_1[20] <= conv1_result[5][2+cnt1][0+cnt2];\
                    producted_1[21] <= conv1_result[5][2+cnt1][1+cnt2];\
                    producted_1[22] <= conv1_result[5][2+cnt1][2+cnt2];\
                    producted_1[23] <= conv1_result[5][2+cnt1][3+cnt2];\
                    producted_1[24] <= conv1_result[5][2+cnt1][4+cnt2];\
                    producted_1[25] <= conv1_result[5][2+cnt1][5+cnt2];\
                    producted_1[26] <= conv1_result[5][2+cnt1][6+cnt2];\
                    producted_1[27] <= conv1_result[5][2+cnt1][7+cnt2];\
                    producted_1[28] <= conv1_result[5][2+cnt1][8+cnt2];\
                    producted_1[29] <= conv1_result[5][2+cnt1][9+cnt2];\
                    producted_1[30] <= conv1_result[5][3+cnt1][0+cnt2];\
                    producted_1[31] <= conv1_result[5][3+cnt1][1+cnt2];\
                    producted_1[32] <= conv1_result[5][3+cnt1][2+cnt2];\
                    producted_1[33] <= conv1_result[5][3+cnt1][3+cnt2];\
                    producted_1[34] <= conv1_result[5][3+cnt1][4+cnt2];\
                    producted_1[35] <= conv1_result[5][3+cnt1][5+cnt2];\
                    producted_1[36] <= conv1_result[5][3+cnt1][6+cnt2];\
                    producted_1[37] <= conv1_result[5][3+cnt1][7+cnt2];\
                    producted_1[38] <= conv1_result[5][3+cnt1][8+cnt2];\
                    producted_1[39] <= conv1_result[5][3+cnt1][9+cnt2];\
                    producted_1[40] <= conv1_result[5][4+cnt1][0+cnt2];\
                    producted_1[41] <= conv1_result[5][4+cnt1][1+cnt2];\
                    producted_1[42] <= conv1_result[5][4+cnt1][2+cnt2];\
                    producted_1[43] <= conv1_result[5][4+cnt1][3+cnt2];\
                    producted_1[44] <= conv1_result[5][4+cnt1][4+cnt2];\
                    producted_1[45] <= conv1_result[5][4+cnt1][5+cnt2];\
                    producted_1[46] <= conv1_result[5][4+cnt1][6+cnt2];\
                    producted_1[47] <= conv1_result[5][4+cnt1][7+cnt2];\
                    producted_1[48] <= conv1_result[5][4+cnt1][8+cnt2];\
                    producted_1[49] <= conv1_result[5][4+cnt1][9+cnt2];\
                    producted_1[50] <= conv1_result[5][5+cnt1][0+cnt2];\
                    producted_1[51] <= conv1_result[5][5+cnt1][1+cnt2];\
                    producted_1[52] <= conv1_result[5][5+cnt1][2+cnt2];\
                    producted_1[53] <= conv1_result[5][5+cnt1][3+cnt2];\
                    producted_1[54] <= conv1_result[5][5+cnt1][4+cnt2];\
                    producted_1[55] <= conv1_result[5][5+cnt1][5+cnt2];\
                    producted_1[56] <= conv1_result[5][5+cnt1][6+cnt2];\
                    producted_1[57] <= conv1_result[5][5+cnt1][7+cnt2];\
                    producted_1[58] <= conv1_result[5][5+cnt1][8+cnt2];\
                    producted_1[59] <= conv1_result[5][5+cnt1][9+cnt2];\
                    producted_1[60] <= conv1_result[5][6+cnt1][0+cnt2];\
                    producted_1[61] <= conv1_result[5][6+cnt1][1+cnt2];\
                    producted_1[62] <= conv1_result[5][6+cnt1][2+cnt2];\
                    producted_1[63] <= conv1_result[5][6+cnt1][3+cnt2];\
                    producted_1[64] <= conv1_result[5][6+cnt1][4+cnt2];\
                    producted_1[65] <= conv1_result[5][6+cnt1][5+cnt2];\
                    producted_1[66] <= conv1_result[5][6+cnt1][6+cnt2];\
                    producted_1[67] <= conv1_result[5][6+cnt1][7+cnt2];\
                    producted_1[68] <= conv1_result[5][6+cnt1][8+cnt2];\
                    producted_1[69] <= conv1_result[5][6+cnt1][9+cnt2];\
                    producted_1[70] <= conv1_result[5][7+cnt1][0+cnt2];\
                    producted_1[71] <= conv1_result[5][7+cnt1][1+cnt2];\
                    producted_1[72] <= conv1_result[5][7+cnt1][2+cnt2];\
                    producted_1[73] <= conv1_result[5][7+cnt1][3+cnt2];\
                    producted_1[74] <= conv1_result[5][7+cnt1][4+cnt2];\
                    producted_1[75] <= conv1_result[5][7+cnt1][5+cnt2];\
                    producted_1[76] <= conv1_result[5][7+cnt1][6+cnt2];\
                    producted_1[77] <= conv1_result[5][7+cnt1][7+cnt2];\
                    producted_1[78] <= conv1_result[5][7+cnt1][8+cnt2];\
                    producted_1[79] <= conv1_result[5][7+cnt1][9+cnt2];\
                    producted_1[80] <= conv1_result[5][8+cnt1][0+cnt2];\
                    producted_1[81] <= conv1_result[5][8+cnt1][1+cnt2];\
                    producted_1[82] <= conv1_result[5][8+cnt1][2+cnt2];\
                    producted_1[83] <= conv1_result[5][8+cnt1][3+cnt2];\
                    producted_1[84] <= conv1_result[5][8+cnt1][4+cnt2];\
                    producted_1[85] <= conv1_result[5][8+cnt1][5+cnt2];\
                    producted_1[86] <= conv1_result[5][8+cnt1][6+cnt2];\
                    producted_1[87] <= conv1_result[5][8+cnt1][7+cnt2];\
                    producted_1[88] <= conv1_result[5][8+cnt1][8+cnt2];\
                    producted_1[89] <= conv1_result[5][8+cnt1][9+cnt2];\
                    producted_1[90] <= conv1_result[5][9+cnt1][0+cnt2];\
                    producted_1[91] <= conv1_result[5][9+cnt1][1+cnt2];\
                    producted_1[92] <= conv1_result[5][9+cnt1][2+cnt2];\
                    producted_1[93] <= conv1_result[5][9+cnt1][3+cnt2];\
                    producted_1[94] <= conv1_result[5][9+cnt1][4+cnt2];\
                    producted_1[95] <= conv1_result[5][9+cnt1][5+cnt2];\
                    producted_1[96] <= conv1_result[5][9+cnt1][6+cnt2];\
                    producted_1[97] <= conv1_result[5][9+cnt1][7+cnt2];\
                    producted_1[98] <= conv1_result[5][9+cnt1][8+cnt2];\
                    producted_1[99] <= conv1_result[5][9+cnt1][9+cnt2];\
					producted_1[100] <= 18'd0;\
					producted_1[101] <= 18'd0;\
					producted_1[102] <= 18'd0;\
					producted_1[103] <= 18'd0;\
					producted_1[104] <= 18'd0;\
					producted_1[105] <= 18'd0;\
					producted_1[106] <= 18'd0;\
					producted_1[107] <= 18'd0;\
					producted_1[108] <= 18'd0;\
					producted_1[109] <= 18'd0;\
					producted_1[110] <= 18'd0;\
					producted_1[111] <= 18'd0;\
                end\
            end\
            LINEAR1  :begin\
				if(cnt1<8'd150) begin\
					producted_1[100] <= conv2_result[cnt1];\
					producted_1[101] <= conv2_result[cnt1];\
					producted_1[102] <= conv2_result[cnt1];\
					producted_1[103] <= conv2_result[cnt1];\
					producted_1[104] <= conv2_result[cnt1];\
					producted_1[105] <= conv2_result[cnt1];\
					producted_1[106] <= conv2_result[cnt1];\
					producted_1[107] <= conv2_result[cnt1];\
					producted_1[108] <= conv2_result[cnt1];\
					producted_1[109] <= conv2_result[cnt1];\
					producted_1[110] <= conv2_result[cnt1];\
					producted_1[111] <= conv2_result[cnt1];\
				end\
			end\
            LINEAR2  :begin\
				if(cnt2<8'd12) begin\
					producted_1[100] <= cache[cnt2+8'd100];\
					producted_1[101] <= cache[cnt2+8'd100];\
					producted_1[102] <= cache[cnt2+8'd100];\
					producted_1[103] <= cache[cnt2+8'd100];\
					producted_1[104] <= cache[cnt2+8'd100];\
					producted_1[105] <= cache[cnt2+8'd100];\
					producted_1[106] <= cache[cnt2+8'd100];\
					producted_1[107] <= cache[cnt2+8'd100];\
					producted_1[108] <= cache[cnt2+8'd100];\
					producted_1[109] <= cache[cnt2+8'd100];\
					producted_1[110] <= 18'd0;\
					producted_1[111] <= 18'd0;\
				end\
			end\
			COMPARE	 :;\
            COMPLETE :;\
            default: begin\
				producted_1[0] <= 18'd0;\
				producted_1[1] <= 18'd0;\
				producted_1[2] <= 18'd0;\
				producted_1[3] <= 18'd0;\
				producted_1[4] <= 18'd0;\
				producted_1[5] <= 18'd0;\
				producted_1[6] <= 18'd0;\
				producted_1[7] <= 18'd0;\
				producted_1[8] <= 18'd0;\
				producted_1[9] <= 18'd0;\
				producted_1[10] <= 18'd0;\
				producted_1[11] <= 18'd0;\
				producted_1[12] <= 18'd0;\
				producted_1[13] <= 18'd0;\
				producted_1[14] <= 18'd0;\
				producted_1[15] <= 18'd0;\
				producted_1[16] <= 18'd0;\
				producted_1[17] <= 18'd0;\
				producted_1[18] <= 18'd0;\
				producted_1[19] <= 18'd0;\
				producted_1[20] <= 18'd0;\
				producted_1[21] <= 18'd0;\
				producted_1[22] <= 18'd0;\
				producted_1[23] <= 18'd0;\
				producted_1[24] <= 18'd0;\
				producted_1[25] <= 18'd0;\
				producted_1[26] <= 18'd0;\
				producted_1[27] <= 18'd0;\
				producted_1[28] <= 18'd0;\
				producted_1[29] <= 18'd0;\
				producted_1[30] <= 18'd0;\
				producted_1[31] <= 18'd0;\
				producted_1[32] <= 18'd0;\
				producted_1[33] <= 18'd0;\
				producted_1[34] <= 18'd0;\
				producted_1[35] <= 18'd0;\
				producted_1[36] <= 18'd0;\
				producted_1[37] <= 18'd0;\
				producted_1[38] <= 18'd0;\
				producted_1[39] <= 18'd0;\
				producted_1[40] <= 18'd0;\
				producted_1[41] <= 18'd0;\
				producted_1[42] <= 18'd0;\
				producted_1[43] <= 18'd0;\
				producted_1[44] <= 18'd0;\
				producted_1[45] <= 18'd0;\
				producted_1[46] <= 18'd0;\
				producted_1[47] <= 18'd0;\
				producted_1[48] <= 18'd0;\
				producted_1[49] <= 18'd0;\
				producted_1[50] <= 18'd0;\
				producted_1[51] <= 18'd0;\
				producted_1[52] <= 18'd0;\
				producted_1[53] <= 18'd0;\
				producted_1[54] <= 18'd0;\
				producted_1[55] <= 18'd0;\
				producted_1[56] <= 18'd0;\
				producted_1[57] <= 18'd0;\
				producted_1[58] <= 18'd0;\
				producted_1[59] <= 18'd0;\
				producted_1[60] <= 18'd0;\
				producted_1[61] <= 18'd0;\
				producted_1[62] <= 18'd0;\
				producted_1[63] <= 18'd0;\
				producted_1[64] <= 18'd0;\
				producted_1[65] <= 18'd0;\
				producted_1[66] <= 18'd0;\
				producted_1[67] <= 18'd0;\
				producted_1[68] <= 18'd0;\
				producted_1[69] <= 18'd0;\
				producted_1[70] <= 18'd0;\
				producted_1[71] <= 18'd0;\
				producted_1[72] <= 18'd0;\
				producted_1[73] <= 18'd0;\
				producted_1[74] <= 18'd0;\
				producted_1[75] <= 18'd0;\
				producted_1[76] <= 18'd0;\
				producted_1[77] <= 18'd0;\
				producted_1[78] <= 18'd0;\
				producted_1[79] <= 18'd0;\
				producted_1[80] <= 18'd0;\
				producted_1[81] <= 18'd0;\
				producted_1[82] <= 18'd0;\
				producted_1[83] <= 18'd0;\
				producted_1[84] <= 18'd0;\
				producted_1[85] <= 18'd0;\
				producted_1[86] <= 18'd0;\
				producted_1[87] <= 18'd0;\
				producted_1[88] <= 18'd0;\
				producted_1[89] <= 18'd0;\
				producted_1[90] <= 18'd0;\
				producted_1[91] <= 18'd0;\
				producted_1[92] <= 18'd0;\
				producted_1[93] <= 18'd0;\
				producted_1[94] <= 18'd0;\
				producted_1[95] <= 18'd0;\
				producted_1[96] <= 18'd0;\
				producted_1[97] <= 18'd0;\
				producted_1[98] <= 18'd0;\
				producted_1[99] <= 18'd0;\
				producted_1[100] <= 18'd0;\
				producted_1[101] <= 18'd0;\
				producted_1[102] <= 18'd0;\
				producted_1[103] <= 18'd0;\
				producted_1[104] <= 18'd0;\
				producted_1[105] <= 18'd0;\
				producted_1[106] <= 18'd0;\
				producted_1[107] <= 18'd0;\
				producted_1[108] <= 18'd0;\
				producted_1[109] <= 18'd0;\
				producted_1[110] <= 18'd0;\
				producted_1[111] <= 18'd0;\
			end\
        endcase\
    end\
end\
always@(posedge clk or negedge rst_n) begin\
    if(!rst_n) begin\
		producted_2[0] <= 18'd0;\
		producted_2[1] <= 18'd0;\
		producted_2[2] <= 18'd0;\
		producted_2[3] <= 18'd0;\
		producted_2[4] <= 18'd0;\
		producted_2[5] <= 18'd0;\
		producted_2[6] <= 18'd0;\
		producted_2[7] <= 18'd0;\
		producted_2[8] <= 18'd0;\
		producted_2[9] <= 18'd0;\
		producted_2[10] <= 18'd0;\
		producted_2[11] <= 18'd0;\
		producted_2[12] <= 18'd0;\
		producted_2[13] <= 18'd0;\
		producted_2[14] <= 18'd0;\
		producted_2[15] <= 18'd0;\
		producted_2[16] <= 18'd0;\
		producted_2[17] <= 18'd0;\
		producted_2[18] <= 18'd0;\
		producted_2[19] <= 18'd0;\
		producted_2[20] <= 18'd0;\
		producted_2[21] <= 18'd0;\
		producted_2[22] <= 18'd0;\
		producted_2[23] <= 18'd0;\
		producted_2[24] <= 18'd0;\
		producted_2[25] <= 18'd0;\
		producted_2[26] <= 18'd0;\
		producted_2[27] <= 18'd0;\
		producted_2[28] <= 18'd0;\
		producted_2[29] <= 18'd0;\
		producted_2[30] <= 18'd0;\
		producted_2[31] <= 18'd0;\
		producted_2[32] <= 18'd0;\
		producted_2[33] <= 18'd0;\
		producted_2[34] <= 18'd0;\
		producted_2[35] <= 18'd0;\
		producted_2[36] <= 18'd0;\
		producted_2[37] <= 18'd0;\
		producted_2[38] <= 18'd0;\
		producted_2[39] <= 18'd0;\
		producted_2[40] <= 18'd0;\
		producted_2[41] <= 18'd0;\
		producted_2[42] <= 18'd0;\
		producted_2[43] <= 18'd0;\
		producted_2[44] <= 18'd0;\
		producted_2[45] <= 18'd0;\
		producted_2[46] <= 18'd0;\
		producted_2[47] <= 18'd0;\
		producted_2[48] <= 18'd0;\
		producted_2[49] <= 18'd0;\
		producted_2[50] <= 18'd0;\
		producted_2[51] <= 18'd0;\
		producted_2[52] <= 18'd0;\
		producted_2[53] <= 18'd0;\
		producted_2[54] <= 18'd0;\
		producted_2[55] <= 18'd0;\
		producted_2[56] <= 18'd0;\
		producted_2[57] <= 18'd0;\
		producted_2[58] <= 18'd0;\
		producted_2[59] <= 18'd0;\
		producted_2[60] <= 18'd0;\
		producted_2[61] <= 18'd0;\
		producted_2[62] <= 18'd0;\
		producted_2[63] <= 18'd0;\
		producted_2[64] <= 18'd0;\
		producted_2[65] <= 18'd0;\
		producted_2[66] <= 18'd0;\
		producted_2[67] <= 18'd0;\
		producted_2[68] <= 18'd0;\
		producted_2[69] <= 18'd0;\
		producted_2[70] <= 18'd0;\
		producted_2[71] <= 18'd0;\
		producted_2[72] <= 18'd0;\
		producted_2[73] <= 18'd0;\
		producted_2[74] <= 18'd0;\
		producted_2[75] <= 18'd0;\
		producted_2[76] <= 18'd0;\
		producted_2[77] <= 18'd0;\
		producted_2[78] <= 18'd0;\
		producted_2[79] <= 18'd0;\
		producted_2[80] <= 18'd0;\
		producted_2[81] <= 18'd0;\
		producted_2[82] <= 18'd0;\
		producted_2[83] <= 18'd0;\
		producted_2[84] <= 18'd0;\
		producted_2[85] <= 18'd0;\
		producted_2[86] <= 18'd0;\
		producted_2[87] <= 18'd0;\
		producted_2[88] <= 18'd0;\
		producted_2[89] <= 18'd0;\
		producted_2[90] <= 18'd0;\
		producted_2[91] <= 18'd0;\
		producted_2[92] <= 18'd0;\
		producted_2[93] <= 18'd0;\
		producted_2[94] <= 18'd0;\
		producted_2[95] <= 18'd0;\
		producted_2[96] <= 18'd0;\
		producted_2[97] <= 18'd0;\
		producted_2[98] <= 18'd0;\
		producted_2[99] <= 18'd0;\
		producted_2[100] <= 18'd0;\
		producted_2[101] <= 18'd0;\
		producted_2[102] <= 18'd0;\
		producted_2[103] <= 18'd0;\
		producted_2[104] <= 18'd0;\
		producted_2[105] <= 18'd0;\
		producted_2[106] <= 18'd0;\
		producted_2[107] <= 18'd0;\
		producted_2[108] <= 18'd0;\
		producted_2[109] <= 18'd0;\
		producted_2[110] <= 18'd0;\
		producted_2[111] <= 18'd0;\
    end\
    else begin\
        case(state)\
            IDLE     :;\
            INPUT    :;\
            CONV1_1_1,CONV1_1_2,CONV1_1_3,CONV1_1_4,CONV1_1_5,CONV1_1_6,CONV1_1_7:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_2[0] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[1] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[2] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[3] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[4] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[5] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[6] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[7] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[8] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[9] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[10] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[11] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[12] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[13] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[14] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[15] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[16] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[17] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[18] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[19] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[20] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[21] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[22] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[23] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[24] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[25] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[26] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[27] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[28] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[29] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[30] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[31] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[32] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[33] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[34] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[35] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[36] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[37] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[38] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[39] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[40] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[41] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[42] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[43] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[44] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[45] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[46] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[47] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[48] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[49] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[50] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[51] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[52] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[53] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[54] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[55] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[56] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[57] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[58] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[59] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[60] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[61] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[62] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[63] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[64] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[65] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[66] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[67] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[68] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[69] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[70] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[71] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[72] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[73] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[74] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[75] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[76] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[77] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[78] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[79] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[80] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[81] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[82] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[83] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[84] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[85] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[86] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[87] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[88] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[89] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[90] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[91] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[92] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[93] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[94] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[95] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[96] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[97] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[98] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[99] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[100] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[101] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[102] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[103] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[104] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[105] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[106] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[107] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[108] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[109] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[110] <= conv1_weight_array[0][cnt1][cnt2];\
					producted_2[111] <= conv1_weight_array[0][cnt1][cnt2];\
                end\
            end\
            CONV1_2_1,CONV1_2_2,CONV1_2_3,CONV1_2_4,CONV1_2_5,CONV1_2_6,CONV1_2_7:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_2[0] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[1] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[2] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[3] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[4] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[5] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[6] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[7] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[8] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[9] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[10] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[11] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[12] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[13] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[14] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[15] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[16] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[17] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[18] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[19] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[20] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[21] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[22] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[23] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[24] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[25] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[26] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[27] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[28] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[29] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[30] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[31] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[32] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[33] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[34] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[35] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[36] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[37] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[38] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[39] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[40] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[41] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[42] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[43] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[44] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[45] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[46] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[47] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[48] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[49] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[50] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[51] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[52] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[53] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[54] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[55] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[56] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[57] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[58] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[59] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[60] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[61] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[62] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[63] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[64] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[65] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[66] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[67] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[68] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[69] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[70] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[71] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[72] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[73] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[74] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[75] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[76] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[77] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[78] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[79] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[80] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[81] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[82] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[83] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[84] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[85] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[86] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[87] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[88] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[89] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[90] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[91] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[92] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[93] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[94] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[95] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[96] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[97] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[98] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[99] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[100] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[101] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[102] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[103] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[104] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[105] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[106] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[107] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[108] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[109] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[110] <= conv1_weight_array[1][cnt1][cnt2];\
					producted_2[111] <= conv1_weight_array[1][cnt1][cnt2];\
                end\
            end\
            CONV1_3_1,CONV1_3_2,CONV1_3_3,CONV1_3_4,CONV1_3_5,CONV1_3_6,CONV1_3_7:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_2[0] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[1] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[2] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[3] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[4] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[5] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[6] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[7] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[8] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[9] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[10] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[11] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[12] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[13] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[14] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[15] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[16] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[17] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[18] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[19] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[20] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[21] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[22] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[23] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[24] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[25] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[26] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[27] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[28] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[29] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[30] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[31] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[32] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[33] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[34] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[35] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[36] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[37] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[38] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[39] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[40] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[41] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[42] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[43] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[44] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[45] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[46] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[47] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[48] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[49] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[50] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[51] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[52] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[53] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[54] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[55] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[56] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[57] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[58] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[59] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[60] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[61] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[62] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[63] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[64] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[65] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[66] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[67] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[68] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[69] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[70] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[71] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[72] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[73] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[74] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[75] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[76] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[77] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[78] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[79] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[80] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[81] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[82] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[83] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[84] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[85] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[86] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[87] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[88] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[89] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[90] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[91] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[92] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[93] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[94] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[95] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[96] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[97] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[98] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[99] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[100] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[101] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[102] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[103] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[104] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[105] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[106] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[107] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[108] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[109] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[110] <= conv1_weight_array[2][cnt1][cnt2];\
					producted_2[111] <= conv1_weight_array[2][cnt1][cnt2];\
                end\
            end\
            CONV1_4_1,CONV1_4_2,CONV1_4_3,CONV1_4_4,CONV1_4_5,CONV1_4_6,CONV1_4_7:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_2[0] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[1] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[2] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[3] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[4] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[5] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[6] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[7] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[8] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[9] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[10] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[11] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[12] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[13] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[14] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[15] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[16] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[17] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[18] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[19] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[20] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[21] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[22] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[23] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[24] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[25] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[26] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[27] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[28] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[29] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[30] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[31] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[32] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[33] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[34] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[35] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[36] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[37] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[38] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[39] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[40] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[41] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[42] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[43] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[44] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[45] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[46] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[47] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[48] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[49] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[50] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[51] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[52] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[53] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[54] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[55] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[56] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[57] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[58] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[59] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[60] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[61] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[62] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[63] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[64] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[65] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[66] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[67] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[68] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[69] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[70] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[71] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[72] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[73] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[74] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[75] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[76] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[77] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[78] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[79] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[80] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[81] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[82] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[83] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[84] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[85] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[86] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[87] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[88] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[89] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[90] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[91] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[92] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[93] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[94] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[95] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[96] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[97] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[98] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[99] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[100] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[101] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[102] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[103] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[104] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[105] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[106] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[107] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[108] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[109] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[110] <= conv1_weight_array[3][cnt1][cnt2];\
					producted_2[111] <= conv1_weight_array[3][cnt1][cnt2];\
                end\
            end\
            CONV1_5_1,CONV1_5_2,CONV1_5_3,CONV1_5_4,CONV1_5_5,CONV1_5_6,CONV1_5_7:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_2[0] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[1] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[2] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[3] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[4] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[5] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[6] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[7] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[8] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[9] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[10] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[11] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[12] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[13] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[14] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[15] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[16] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[17] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[18] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[19] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[20] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[21] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[22] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[23] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[24] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[25] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[26] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[27] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[28] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[29] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[30] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[31] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[32] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[33] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[34] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[35] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[36] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[37] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[38] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[39] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[40] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[41] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[42] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[43] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[44] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[45] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[46] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[47] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[48] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[49] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[50] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[51] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[52] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[53] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[54] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[55] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[56] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[57] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[58] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[59] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[60] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[61] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[62] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[63] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[64] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[65] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[66] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[67] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[68] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[69] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[70] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[71] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[72] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[73] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[74] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[75] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[76] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[77] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[78] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[79] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[80] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[81] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[82] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[83] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[84] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[85] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[86] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[87] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[88] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[89] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[90] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[91] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[92] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[93] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[94] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[95] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[96] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[97] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[98] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[99] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[100] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[101] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[102] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[103] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[104] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[105] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[106] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[107] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[108] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[109] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[110] <= conv1_weight_array[4][cnt1][cnt2];\
					producted_2[111] <= conv1_weight_array[4][cnt1][cnt2];\
                end\
            end\
            CONV1_6_1,CONV1_6_2,CONV1_6_3,CONV1_6_4,CONV1_6_5,CONV1_6_6,CONV1_6_7:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
					producted_2[0] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[1] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[2] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[3] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[4] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[5] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[6] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[7] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[8] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[9] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[10] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[11] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[12] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[13] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[14] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[15] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[16] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[17] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[18] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[19] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[20] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[21] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[22] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[23] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[24] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[25] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[26] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[27] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[28] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[29] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[30] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[31] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[32] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[33] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[34] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[35] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[36] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[37] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[38] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[39] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[40] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[41] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[42] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[43] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[44] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[45] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[46] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[47] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[48] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[49] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[50] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[51] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[52] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[53] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[54] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[55] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[56] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[57] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[58] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[59] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[60] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[61] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[62] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[63] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[64] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[65] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[66] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[67] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[68] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[69] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[70] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[71] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[72] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[73] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[74] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[75] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[76] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[77] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[78] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[79] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[80] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[81] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[82] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[83] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[84] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[85] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[86] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[87] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[88] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[89] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[90] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[91] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[92] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[93] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[94] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[95] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[96] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[97] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[98] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[99] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[100] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[101] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[102] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[103] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[104] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[105] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[106] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[107] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[108] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[109] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[110] <= conv1_weight_array[5][cnt1][cnt2];\
					producted_2[111] <= conv1_weight_array[5][cnt1][cnt2];\
                end\
            end\
            CONV2_1_1:begin\
				producted_2[ 0] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[0][0][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_1_2:begin\
				producted_2[ 0] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[0][1][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_1_3:begin\
				producted_2[ 0] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[0][2][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_1_4:begin\
				producted_2[ 0] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[0][3][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_1_5:begin\
				producted_2[ 0] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[0][4][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_1_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_2[ 0] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 1] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 2] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 3] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 4] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 5] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 6] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 7] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 8] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[ 9] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[10] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[11] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[12] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[13] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[14] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[15] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[16] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[17] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[18] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[19] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[20] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[21] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[22] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[23] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[24] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[25] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[26] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[27] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[28] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[29] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[30] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[31] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[32] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[33] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[34] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[35] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[36] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[37] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[38] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[39] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[40] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[41] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[42] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[43] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[44] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[45] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[46] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[47] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[48] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[49] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[50] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[51] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[52] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[53] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[54] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[55] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[56] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[57] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[58] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[59] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[60] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[61] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[62] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[63] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[64] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[65] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[66] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[67] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[68] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[69] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[70] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[71] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[72] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[73] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[74] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[75] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[76] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[77] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[78] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[79] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[80] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[81] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[82] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[83] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[84] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[85] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[86] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[87] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[88] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[89] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[90] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[91] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[92] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[93] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[94] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[95] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[96] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[97] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[98] <= conv2_weight_array[0][5][cnt1][cnt2];\
                    producted_2[99] <= conv2_weight_array[0][5][cnt1][cnt2];\
					producted_2[100] <= 18'd0;\
					producted_2[101] <= 18'd0;\
					producted_2[102] <= 18'd0;\
					producted_2[103] <= 18'd0;\
					producted_2[104] <= 18'd0;\
					producted_2[105] <= 18'd0;\
					producted_2[106] <= 18'd0;\
					producted_2[107] <= 18'd0;\
					producted_2[108] <= 18'd0;\
					producted_2[109] <= 18'd0;\
					producted_2[110] <= 18'd0;\
					producted_2[111] <= 18'd0;\
                end\
            end\
            CONV2_2_1:begin\
				producted_2[ 0] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[1][0][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_2_2:begin\
				producted_2[ 0] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[1][1][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_2_3:begin\
				producted_2[ 0] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[1][2][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_2_4:begin\
				producted_2[ 0] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[1][3][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_2_5:begin\
				producted_2[ 0] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[1][4][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_2_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_2[ 0] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 1] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 2] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 3] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 4] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 5] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 6] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 7] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 8] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[ 9] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[10] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[11] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[12] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[13] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[14] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[15] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[16] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[17] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[18] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[19] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[20] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[21] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[22] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[23] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[24] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[25] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[26] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[27] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[28] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[29] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[30] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[31] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[32] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[33] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[34] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[35] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[36] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[37] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[38] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[39] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[40] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[41] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[42] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[43] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[44] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[45] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[46] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[47] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[48] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[49] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[50] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[51] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[52] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[53] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[54] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[55] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[56] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[57] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[58] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[59] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[60] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[61] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[62] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[63] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[64] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[65] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[66] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[67] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[68] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[69] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[70] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[71] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[72] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[73] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[74] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[75] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[76] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[77] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[78] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[79] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[80] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[81] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[82] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[83] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[84] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[85] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[86] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[87] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[88] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[89] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[90] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[91] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[92] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[93] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[94] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[95] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[96] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[97] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[98] <= conv2_weight_array[1][5][cnt1][cnt2];\
                    producted_2[99] <= conv2_weight_array[1][5][cnt1][cnt2];\
					producted_2[100] <= 18'd0;\
					producted_2[101] <= 18'd0;\
					producted_2[102] <= 18'd0;\
					producted_2[103] <= 18'd0;\
					producted_2[104] <= 18'd0;\
					producted_2[105] <= 18'd0;\
					producted_2[106] <= 18'd0;\
					producted_2[107] <= 18'd0;\
					producted_2[108] <= 18'd0;\
					producted_2[109] <= 18'd0;\
					producted_2[110] <= 18'd0;\
					producted_2[111] <= 18'd0;\
                end\
            end\
            CONV2_3_1:begin\
				producted_2[ 0] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[2][0][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_3_2:begin\
				producted_2[ 0] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[2][1][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
			end\
            CONV2_3_3:begin\
				producted_2[ 0] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[2][2][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_3_4:begin\
				producted_2[ 0] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[2][3][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_3_5:begin\
				producted_2[ 0] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[2][4][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_3_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_2[ 0] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 1] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 2] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 3] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 4] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 5] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 6] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 7] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 8] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[ 9] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[10] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[11] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[12] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[13] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[14] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[15] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[16] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[17] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[18] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[19] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[20] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[21] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[22] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[23] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[24] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[25] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[26] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[27] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[28] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[29] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[30] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[31] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[32] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[33] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[34] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[35] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[36] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[37] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[38] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[39] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[40] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[41] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[42] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[43] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[44] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[45] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[46] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[47] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[48] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[49] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[50] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[51] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[52] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[53] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[54] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[55] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[56] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[57] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[58] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[59] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[60] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[61] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[62] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[63] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[64] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[65] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[66] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[67] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[68] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[69] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[70] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[71] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[72] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[73] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[74] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[75] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[76] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[77] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[78] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[79] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[80] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[81] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[82] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[83] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[84] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[85] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[86] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[87] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[88] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[89] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[90] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[91] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[92] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[93] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[94] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[95] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[96] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[97] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[98] <= conv2_weight_array[2][5][cnt1][cnt2];\
                    producted_2[99] <= conv2_weight_array[2][5][cnt1][cnt2];\
					producted_2[100] <= 18'd0;\
					producted_2[101] <= 18'd0;\
					producted_2[102] <= 18'd0;\
					producted_2[103] <= 18'd0;\
					producted_2[104] <= 18'd0;\
					producted_2[105] <= 18'd0;\
					producted_2[106] <= 18'd0;\
					producted_2[107] <= 18'd0;\
					producted_2[108] <= 18'd0;\
					producted_2[109] <= 18'd0;\
					producted_2[110] <= 18'd0;\
					producted_2[111] <= 18'd0;\
                end\
            end\
            CONV2_4_1:begin\
				producted_2[ 0] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[3][0][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_4_2:begin\
				producted_2[ 0] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[3][1][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_4_3:begin\
				producted_2[ 0] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[3][2][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_4_4:begin\
				producted_2[ 0] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[3][3][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_4_5:begin\
				producted_2[ 0] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[3][4][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_4_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_2[ 0] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 1] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 2] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 3] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 4] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 5] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 6] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 7] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 8] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[ 9] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[10] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[11] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[12] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[13] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[14] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[15] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[16] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[17] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[18] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[19] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[20] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[21] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[22] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[23] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[24] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[25] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[26] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[27] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[28] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[29] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[30] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[31] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[32] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[33] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[34] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[35] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[36] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[37] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[38] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[39] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[40] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[41] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[42] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[43] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[44] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[45] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[46] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[47] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[48] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[49] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[50] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[51] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[52] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[53] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[54] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[55] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[56] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[57] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[58] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[59] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[60] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[61] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[62] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[63] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[64] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[65] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[66] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[67] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[68] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[69] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[70] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[71] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[72] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[73] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[74] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[75] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[76] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[77] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[78] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[79] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[80] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[81] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[82] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[83] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[84] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[85] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[86] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[87] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[88] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[89] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[90] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[91] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[92] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[93] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[94] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[95] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[96] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[97] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[98] <= conv2_weight_array[3][5][cnt1][cnt2];\
                    producted_2[99] <= conv2_weight_array[3][5][cnt1][cnt2];\
					producted_2[100] <= 18'd0;\
					producted_2[101] <= 18'd0;\
					producted_2[102] <= 18'd0;\
					producted_2[103] <= 18'd0;\
					producted_2[104] <= 18'd0;\
					producted_2[105] <= 18'd0;\
					producted_2[106] <= 18'd0;\
					producted_2[107] <= 18'd0;\
					producted_2[108] <= 18'd0;\
					producted_2[109] <= 18'd0;\
					producted_2[110] <= 18'd0;\
					producted_2[111] <= 18'd0;\
                end\
            end\
            CONV2_5_1:begin\
				producted_2[ 0] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[4][0][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_5_2:begin\
				producted_2[ 0] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[4][1][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_5_3:begin\
				producted_2[ 0] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[4][2][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_5_4:begin\
				producted_2[ 0] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[4][3][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_5_5:begin\
				producted_2[ 0] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[4][4][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_5_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_2[ 0] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 1] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 2] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 3] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 4] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 5] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 6] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 7] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 8] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[ 9] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[10] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[11] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[12] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[13] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[14] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[15] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[16] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[17] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[18] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[19] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[20] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[21] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[22] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[23] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[24] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[25] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[26] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[27] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[28] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[29] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[30] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[31] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[32] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[33] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[34] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[35] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[36] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[37] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[38] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[39] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[40] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[41] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[42] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[43] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[44] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[45] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[46] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[47] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[48] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[49] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[50] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[51] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[52] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[53] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[54] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[55] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[56] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[57] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[58] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[59] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[60] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[61] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[62] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[63] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[64] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[65] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[66] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[67] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[68] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[69] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[70] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[71] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[72] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[73] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[74] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[75] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[76] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[77] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[78] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[79] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[80] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[81] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[82] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[83] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[84] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[85] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[86] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[87] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[88] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[89] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[90] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[91] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[92] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[93] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[94] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[95] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[96] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[97] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[98] <= conv2_weight_array[4][5][cnt1][cnt2];\
                    producted_2[99] <= conv2_weight_array[4][5][cnt1][cnt2];\
					producted_2[100] <= 18'd0;\
					producted_2[101] <= 18'd0;\
					producted_2[102] <= 18'd0;\
					producted_2[103] <= 18'd0;\
					producted_2[104] <= 18'd0;\
					producted_2[105] <= 18'd0;\
					producted_2[106] <= 18'd0;\
					producted_2[107] <= 18'd0;\
					producted_2[108] <= 18'd0;\
					producted_2[109] <= 18'd0;\
					producted_2[110] <= 18'd0;\
					producted_2[111] <= 18'd0;\
                end\
            end\
            CONV2_6_1:begin\
				producted_2[ 0] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[5][0][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_6_2:begin\
				producted_2[ 0] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[5][1][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_6_3:begin\
				producted_2[ 0] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[5][2][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_6_4:begin\
				producted_2[ 0] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[5][3][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_6_5:begin\
				producted_2[ 0] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 1] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 2] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 3] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 4] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 5] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 6] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 7] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 8] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[ 9] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[10] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[11] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[12] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[13] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[14] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[15] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[16] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[17] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[18] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[19] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[20] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[21] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[22] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[23] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[24] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[25] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[26] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[27] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[28] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[29] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[30] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[31] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[32] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[33] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[34] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[35] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[36] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[37] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[38] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[39] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[40] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[41] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[42] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[43] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[44] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[45] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[46] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[47] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[48] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[49] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[50] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[51] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[52] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[53] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[54] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[55] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[56] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[57] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[58] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[59] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[60] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[61] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[62] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[63] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[64] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[65] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[66] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[67] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[68] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[69] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[70] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[71] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[72] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[73] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[74] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[75] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[76] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[77] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[78] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[79] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[80] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[81] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[82] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[83] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[84] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[85] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[86] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[87] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[88] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[89] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[90] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[91] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[92] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[93] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[94] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[95] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[96] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[97] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[98] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[99] <= conv2_weight_array[5][4][cnt1][cnt2];\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
            end\
            CONV2_6_6:begin\
                if((cnt1<=8'd4)&(cnt2<=8'd4)) begin\
                    producted_2[ 0] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 1] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 2] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 3] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 4] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 5] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 6] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 7] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 8] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[ 9] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[10] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[11] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[12] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[13] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[14] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[15] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[16] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[17] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[18] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[19] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[20] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[21] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[22] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[23] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[24] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[25] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[26] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[27] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[28] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[29] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[30] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[31] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[32] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[33] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[34] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[35] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[36] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[37] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[38] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[39] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[40] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[41] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[42] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[43] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[44] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[45] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[46] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[47] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[48] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[49] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[50] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[51] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[52] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[53] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[54] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[55] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[56] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[57] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[58] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[59] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[60] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[61] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[62] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[63] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[64] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[65] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[66] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[67] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[68] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[69] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[70] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[71] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[72] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[73] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[74] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[75] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[76] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[77] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[78] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[79] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[80] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[81] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[82] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[83] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[84] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[85] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[86] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[87] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[88] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[89] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[90] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[91] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[92] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[93] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[94] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[95] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[96] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[97] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[98] <= conv2_weight_array[5][5][cnt1][cnt2];\
                    producted_2[99] <= conv2_weight_array[5][5][cnt1][cnt2];\
					producted_2[100] <= 18'd0;\
					producted_2[101] <= 18'd0;\
					producted_2[102] <= 18'd0;\
					producted_2[103] <= 18'd0;\
					producted_2[104] <= 18'd0;\
					producted_2[105] <= 18'd0;\
					producted_2[106] <= 18'd0;\
					producted_2[107] <= 18'd0;\
					producted_2[108] <= 18'd0;\
					producted_2[109] <= 18'd0;\
					producted_2[110] <= 18'd0;\
					producted_2[111] <= 18'd0;\
                end\
            end\
            LINEAR1  :begin\
				if(cnt1<8'd150) begin\
					producted_2[0] <= 18'd0;\
                    producted_2[1] <= 18'd0;\
                    producted_2[2] <= 18'd0;\
                    producted_2[3] <= 18'd0;\
                    producted_2[4] <= 18'd0;\
                    producted_2[5] <= 18'd0;\
                    producted_2[6] <= 18'd0;\
                    producted_2[7] <= 18'd0;\
                    producted_2[8] <= 18'd0;\
                    producted_2[9] <= 18'd0;\
                    producted_2[10] <= 18'd0;\
                    producted_2[11] <= 18'd0;\
                    producted_2[12] <= 18'd0;\
                    producted_2[13] <= 18'd0;\
                    producted_2[14] <= 18'd0;\
                    producted_2[15] <= 18'd0;\
                    producted_2[16] <= 18'd0;\
                    producted_2[17] <= 18'd0;\
                    producted_2[18] <= 18'd0;\
                    producted_2[19] <= 18'd0;\
                    producted_2[20] <= 18'd0;\
                    producted_2[21] <= 18'd0;\
                    producted_2[22] <= 18'd0;\
                    producted_2[23] <= 18'd0;\
                    producted_2[24] <= 18'd0;\
                    producted_2[25] <= 18'd0;\
                    producted_2[26] <= 18'd0;\
                    producted_2[27] <= 18'd0;\
                    producted_2[28] <= 18'd0;\
                    producted_2[29] <= 18'd0;\
                    producted_2[30] <= 18'd0;\
                    producted_2[31] <= 18'd0;\
                    producted_2[32] <= 18'd0;\
                    producted_2[33] <= 18'd0;\
                    producted_2[34] <= 18'd0;\
                    producted_2[35] <= 18'd0;\
                    producted_2[36] <= 18'd0;\
                    producted_2[37] <= 18'd0;\
                    producted_2[38] <= 18'd0;\
                    producted_2[39] <= 18'd0;\
                    producted_2[40] <= 18'd0;\
                    producted_2[41] <= 18'd0;\
                    producted_2[42] <= 18'd0;\
                    producted_2[43] <= 18'd0;\
                    producted_2[44] <= 18'd0;\
                    producted_2[45] <= 18'd0;\
                    producted_2[46] <= 18'd0;\
                    producted_2[47] <= 18'd0;\
                    producted_2[48] <= 18'd0;\
                    producted_2[49] <= 18'd0;\
                    producted_2[50] <= 18'd0;\
                    producted_2[51] <= 18'd0;\
                    producted_2[52] <= 18'd0;\
                    producted_2[53] <= 18'd0;\
                    producted_2[54] <= 18'd0;\
                    producted_2[55] <= 18'd0;\
                    producted_2[56] <= 18'd0;\
                    producted_2[57] <= 18'd0;\
                    producted_2[58] <= 18'd0;\
                    producted_2[59] <= 18'd0;\
                    producted_2[60] <= 18'd0;\
                    producted_2[61] <= 18'd0;\
                    producted_2[62] <= 18'd0;\
                    producted_2[63] <= 18'd0;\
                    producted_2[64] <= 18'd0;\
                    producted_2[65] <= 18'd0;\
                    producted_2[66] <= 18'd0;\
                    producted_2[67] <= 18'd0;\
                    producted_2[68] <= 18'd0;\
                    producted_2[69] <= 18'd0;\
                    producted_2[70] <= 18'd0;\
                    producted_2[71] <= 18'd0;\
                    producted_2[72] <= 18'd0;\
                    producted_2[73] <= 18'd0;\
                    producted_2[74] <= 18'd0;\
                    producted_2[75] <= 18'd0;\
                    producted_2[76] <= 18'd0;\
                    producted_2[77] <= 18'd0;\
                    producted_2[78] <= 18'd0;\
                    producted_2[79] <= 18'd0;\
                    producted_2[80] <= 18'd0;\
                    producted_2[81] <= 18'd0;\
                    producted_2[82] <= 18'd0;\
                    producted_2[83] <= 18'd0;\
                    producted_2[84] <= 18'd0;\
                    producted_2[85] <= 18'd0;\
                    producted_2[86] <= 18'd0;\
                    producted_2[87] <= 18'd0;\
                    producted_2[88] <= 18'd0;\
                    producted_2[89] <= 18'd0;\
                    producted_2[90] <= 18'd0;\
                    producted_2[91] <= 18'd0;\
                    producted_2[92] <= 18'd0;\
                    producted_2[93] <= 18'd0;\
                    producted_2[94] <= 18'd0;\
                    producted_2[95] <= 18'd0;\
                    producted_2[96] <= 18'd0;\
                    producted_2[97] <= 18'd0;\
                    producted_2[98] <= 18'd0;\
                    producted_2[99] <= 18'd0;\
					producted_2[100] <= linear1_weight_array[0][cnt1];\
					producted_2[101] <= linear1_weight_array[1][cnt1];\
					producted_2[102] <= linear1_weight_array[2][cnt1];\
					producted_2[103] <= linear1_weight_array[3][cnt1];\
					producted_2[104] <= linear1_weight_array[4][cnt1];\
					producted_2[105] <= linear1_weight_array[5][cnt1];\
					producted_2[106] <= linear1_weight_array[6][cnt1];\
					producted_2[107] <= linear1_weight_array[7][cnt1];\
					producted_2[108] <= linear1_weight_array[8][cnt1];\
					producted_2[109] <= linear1_weight_array[9][cnt1];\
					producted_2[110] <= linear1_weight_array[10][cnt1];\
					producted_2[111] <= linear1_weight_array[11][cnt1];\
				end\
			end\
            LINEAR2  :begin\
				if(cnt2<8'd12) begin\
					producted_2[100] <= linear2_weight_array[0][cnt2];\
					producted_2[101] <= linear2_weight_array[1][cnt2];\
					producted_2[102] <= linear2_weight_array[2][cnt2];\
					producted_2[103] <= linear2_weight_array[3][cnt2];\
					producted_2[104] <= linear2_weight_array[4][cnt2];\
					producted_2[105] <= linear2_weight_array[5][cnt2];\
					producted_2[106] <= linear2_weight_array[6][cnt2];\
					producted_2[107] <= linear2_weight_array[7][cnt2];\
					producted_2[108] <= linear2_weight_array[8][cnt2];\
					producted_2[109] <= linear2_weight_array[9][cnt2];\
				end\
			end\
			COMPARE  :;\
            COMPLETE :;\
            default: begin\
				producted_2[0] <= 18'd0;\
				producted_2[1] <= 18'd0;\
				producted_2[2] <= 18'd0;\
				producted_2[3] <= 18'd0;\
				producted_2[4] <= 18'd0;\
				producted_2[5] <= 18'd0;\
				producted_2[6] <= 18'd0;\
				producted_2[7] <= 18'd0;\
				producted_2[8] <= 18'd0;\
				producted_2[9] <= 18'd0;\
				producted_2[10] <= 18'd0;\
				producted_2[11] <= 18'd0;\
				producted_2[12] <= 18'd0;\
				producted_2[13] <= 18'd0;\
				producted_2[14] <= 18'd0;\
				producted_2[15] <= 18'd0;\
				producted_2[16] <= 18'd0;\
				producted_2[17] <= 18'd0;\
				producted_2[18] <= 18'd0;\
				producted_2[19] <= 18'd0;\
				producted_2[20] <= 18'd0;\
				producted_2[21] <= 18'd0;\
				producted_2[22] <= 18'd0;\
				producted_2[23] <= 18'd0;\
				producted_2[24] <= 18'd0;\
				producted_2[25] <= 18'd0;\
				producted_2[26] <= 18'd0;\
				producted_2[27] <= 18'd0;\
				producted_2[28] <= 18'd0;\
				producted_2[29] <= 18'd0;\
				producted_2[30] <= 18'd0;\
				producted_2[31] <= 18'd0;\
				producted_2[32] <= 18'd0;\
				producted_2[33] <= 18'd0;\
				producted_2[34] <= 18'd0;\
				producted_2[35] <= 18'd0;\
				producted_2[36] <= 18'd0;\
				producted_2[37] <= 18'd0;\
				producted_2[38] <= 18'd0;\
				producted_2[39] <= 18'd0;\
				producted_2[40] <= 18'd0;\
				producted_2[41] <= 18'd0;\
				producted_2[42] <= 18'd0;\
				producted_2[43] <= 18'd0;\
				producted_2[44] <= 18'd0;\
				producted_2[45] <= 18'd0;\
				producted_2[46] <= 18'd0;\
				producted_2[47] <= 18'd0;\
				producted_2[48] <= 18'd0;\
				producted_2[49] <= 18'd0;\
				producted_2[50] <= 18'd0;\
				producted_2[51] <= 18'd0;\
				producted_2[52] <= 18'd0;\
				producted_2[53] <= 18'd0;\
				producted_2[54] <= 18'd0;\
				producted_2[55] <= 18'd0;\
				producted_2[56] <= 18'd0;\
				producted_2[57] <= 18'd0;\
				producted_2[58] <= 18'd0;\
				producted_2[59] <= 18'd0;\
				producted_2[60] <= 18'd0;\
				producted_2[61] <= 18'd0;\
				producted_2[62] <= 18'd0;\
				producted_2[63] <= 18'd0;\
				producted_2[64] <= 18'd0;\
				producted_2[65] <= 18'd0;\
				producted_2[66] <= 18'd0;\
				producted_2[67] <= 18'd0;\
				producted_2[68] <= 18'd0;\
				producted_2[69] <= 18'd0;\
				producted_2[70] <= 18'd0;\
				producted_2[71] <= 18'd0;\
				producted_2[72] <= 18'd0;\
				producted_2[73] <= 18'd0;\
				producted_2[74] <= 18'd0;\
				producted_2[75] <= 18'd0;\
				producted_2[76] <= 18'd0;\
				producted_2[77] <= 18'd0;\
				producted_2[78] <= 18'd0;\
				producted_2[79] <= 18'd0;\
				producted_2[80] <= 18'd0;\
				producted_2[81] <= 18'd0;\
				producted_2[82] <= 18'd0;\
				producted_2[83] <= 18'd0;\
				producted_2[84] <= 18'd0;\
				producted_2[85] <= 18'd0;\
				producted_2[86] <= 18'd0;\
				producted_2[87] <= 18'd0;\
				producted_2[88] <= 18'd0;\
				producted_2[89] <= 18'd0;\
				producted_2[90] <= 18'd0;\
				producted_2[91] <= 18'd0;\
				producted_2[92] <= 18'd0;\
				producted_2[93] <= 18'd0;\
				producted_2[94] <= 18'd0;\
				producted_2[95] <= 18'd0;\
				producted_2[96] <= 18'd0;\
				producted_2[97] <= 18'd0;\
				producted_2[98] <= 18'd0;\
				producted_2[99] <= 18'd0;\
				producted_2[100] <= 18'd0;\
				producted_2[101] <= 18'd0;\
				producted_2[102] <= 18'd0;\
				producted_2[103] <= 18'd0;\
				producted_2[104] <= 18'd0;\
				producted_2[105] <= 18'd0;\
				producted_2[106] <= 18'd0;\
				producted_2[107] <= 18'd0;\
				producted_2[108] <= 18'd0;\
				producted_2[109] <= 18'd0;\
				producted_2[110] <= 18'd0;\
				producted_2[111] <= 18'd0;\
			end\
        endcase\
    end\
end