// //kernel = 0.25
// `define CONV2_WEIGHT \
// reg [0:449] conv2_weight_array [0:5][0:5];\
// always@(posedge clk or negedge rst_n) begin\
//     conv2_weight_array[0][0] <= {25{18'h00100}};\
//     conv2_weight_array[0][1] <= {25{18'h00100}};\
//     conv2_weight_array[0][2] <= {25{18'h00100}};\
//     conv2_weight_array[0][3] <= {25{18'h00100}};\
//     conv2_weight_array[0][4] <= {25{18'h00100}};\
//     conv2_weight_array[0][5] <= {25{18'h00100}};\
//     conv2_weight_array[1][0] <= {25{18'h00100}};\
//     conv2_weight_array[1][1] <= {25{18'h00100}};\
//     conv2_weight_array[1][2] <= {25{18'h00100}};\
//     conv2_weight_array[1][3] <= {25{18'h00100}};\
//     conv2_weight_array[1][4] <= {25{18'h00100}};\
//     conv2_weight_array[1][5] <= {25{18'h00100}};\
//     conv2_weight_array[2][0] <= {25{18'h00100}};\
//     conv2_weight_array[2][1] <= {25{18'h00100}};\
//     conv2_weight_array[2][2] <= {25{18'h00100}};\
//     conv2_weight_array[2][3] <= {25{18'h00100}};\
//     conv2_weight_array[2][4] <= {25{18'h00100}};\
//     conv2_weight_array[2][5] <= {25{18'h00100}};\
//     conv2_weight_array[3][0] <= {25{18'h00100}};\
//     conv2_weight_array[3][1] <= {25{18'h00100}};\
//     conv2_weight_array[3][2] <= {25{18'h00100}};\
//     conv2_weight_array[3][3] <= {25{18'h00100}};\
//     conv2_weight_array[3][4] <= {25{18'h00100}};\
//     conv2_weight_array[3][5] <= {25{18'h00100}};\
//     conv2_weight_array[4][0] <= {25{18'h00100}};\
//     conv2_weight_array[4][1] <= {25{18'h00100}};\
//     conv2_weight_array[4][2] <= {25{18'h00100}};\
//     conv2_weight_array[4][3] <= {25{18'h00100}};\
//     conv2_weight_array[4][4] <= {25{18'h00100}};\
//     conv2_weight_array[4][5] <= {25{18'h00100}};\
//     conv2_weight_array[5][0] <= {25{18'h00100}};\
//     conv2_weight_array[5][1] <= {25{18'h00100}};\
//     conv2_weight_array[5][2] <= {25{18'h00100}};\
//     conv2_weight_array[5][3] <= {25{18'h00100}};\
//     conv2_weight_array[5][4] <= {25{18'h00100}};\
//     conv2_weight_array[5][5] <= {25{18'h00100}};\
// end

`define CONV2_WEIGHT \
reg [0:17] conv2_weight_array [0:5][0:5][0:4][0:4];\
always@(posedge clk) begin\
    conv2_weight_array[0][0][0][0] <= 18'b100000000100111101;\
    conv2_weight_array[0][0][0][1] <= 18'b100000000010011011;\
    conv2_weight_array[0][0][0][2] <= 18'b100000000001101000;\
    conv2_weight_array[0][0][0][3] <= 18'b100000000001110111;\
    conv2_weight_array[0][0][0][4] <= 18'b100000000010000000;\
    conv2_weight_array[0][0][1][0] <= 18'b000000000010001110;\
    conv2_weight_array[0][0][1][1] <= 18'b000000000010101101;\
    conv2_weight_array[0][0][1][2] <= 18'b000000000011111100;\
    conv2_weight_array[0][0][1][3] <= 18'b000000000110001001;\
    conv2_weight_array[0][0][1][4] <= 18'b000000000001100111;\
    conv2_weight_array[0][0][2][0] <= 18'b000000000101000110;\
    conv2_weight_array[0][0][2][1] <= 18'b000000000011110110;\
    conv2_weight_array[0][0][2][2] <= 18'b000000000100010000;\
    conv2_weight_array[0][0][2][3] <= 18'b000000000110101101;\
    conv2_weight_array[0][0][2][4] <= 18'b000000001001010010;\
    conv2_weight_array[0][0][3][0] <= 18'b000000000000110010;\
    conv2_weight_array[0][0][3][1] <= 18'b100000000000001111;\
    conv2_weight_array[0][0][3][2] <= 18'b100000000000010111;\
    conv2_weight_array[0][0][3][3] <= 18'b000000000000100111;\
    conv2_weight_array[0][0][3][4] <= 18'b000000000000110100;\
    conv2_weight_array[0][0][4][0] <= 18'b100000000011100101;\
    conv2_weight_array[0][0][4][1] <= 18'b100000000110111111;\
    conv2_weight_array[0][0][4][2] <= 18'b000000000000111001;\
    conv2_weight_array[0][0][4][3] <= 18'b000000000001001011;\
    conv2_weight_array[0][0][4][4] <= 18'b000000000100100100;\
    conv2_weight_array[0][1][0][0] <= 18'b000000000001100111;\
    conv2_weight_array[0][1][0][1] <= 18'b000000000011001000;\
    conv2_weight_array[0][1][0][2] <= 18'b100000001000000011;\
    conv2_weight_array[0][1][0][3] <= 18'b100000000000100111;\
    conv2_weight_array[0][1][0][4] <= 18'b000000001011011011;\
    conv2_weight_array[0][1][1][0] <= 18'b100000000000000010;\
    conv2_weight_array[0][1][1][1] <= 18'b000000000000110111;\
    conv2_weight_array[0][1][1][2] <= 18'b100000000100111111;\
    conv2_weight_array[0][1][1][3] <= 18'b100000001001011001;\
    conv2_weight_array[0][1][1][4] <= 18'b100000001000110001;\
    conv2_weight_array[0][1][2][0] <= 18'b000000000101000111;\
    conv2_weight_array[0][1][2][1] <= 18'b000000000011000101;\
    conv2_weight_array[0][1][2][2] <= 18'b100000000000011110;\
    conv2_weight_array[0][1][2][3] <= 18'b100000000110000000;\
    conv2_weight_array[0][1][2][4] <= 18'b100000000110100110;\
    conv2_weight_array[0][1][3][0] <= 18'b000000000000111010;\
    conv2_weight_array[0][1][3][1] <= 18'b000000000001100010;\
    conv2_weight_array[0][1][3][2] <= 18'b100000000001001110;\
    conv2_weight_array[0][1][3][3] <= 18'b100000000000100110;\
    conv2_weight_array[0][1][3][4] <= 18'b000000000001001000;\
    conv2_weight_array[0][1][4][0] <= 18'b100000000101101100;\
    conv2_weight_array[0][1][4][1] <= 18'b100000000001000000;\
    conv2_weight_array[0][1][4][2] <= 18'b000000000010111011;\
    conv2_weight_array[0][1][4][3] <= 18'b000000000000110000;\
    conv2_weight_array[0][1][4][4] <= 18'b000000000000010110;\
    conv2_weight_array[0][2][0][0] <= 18'b100000000011111010;\
    conv2_weight_array[0][2][0][1] <= 18'b100000000100111100;\
    conv2_weight_array[0][2][0][2] <= 18'b100000000101100100;\
    conv2_weight_array[0][2][0][3] <= 18'b100000000010010011;\
    conv2_weight_array[0][2][0][4] <= 18'b000000000101111001;\
    conv2_weight_array[0][2][1][0] <= 18'b000000000001011110;\
    conv2_weight_array[0][2][1][1] <= 18'b000000000001011010;\
    conv2_weight_array[0][2][1][2] <= 18'b100000000010000111;\
    conv2_weight_array[0][2][1][3] <= 18'b100000000101101001;\
    conv2_weight_array[0][2][1][4] <= 18'b100000001000010010;\
    conv2_weight_array[0][2][2][0] <= 18'b000000000110001010;\
    conv2_weight_array[0][2][2][1] <= 18'b000000000100011110;\
    conv2_weight_array[0][2][2][2] <= 18'b000000000101100001;\
    conv2_weight_array[0][2][2][3] <= 18'b000000000101011101;\
    conv2_weight_array[0][2][2][4] <= 18'b000000000010111100;\
    conv2_weight_array[0][2][3][0] <= 18'b000000000011011110;\
    conv2_weight_array[0][2][3][1] <= 18'b000000000001010001;\
    conv2_weight_array[0][2][3][2] <= 18'b100000000000100011;\
    conv2_weight_array[0][2][3][3] <= 18'b000000000010001110;\
    conv2_weight_array[0][2][3][4] <= 18'b000000000001001001;\
    conv2_weight_array[0][2][4][0] <= 18'b100000000010100001;\
    conv2_weight_array[0][2][4][1] <= 18'b100000000001011010;\
    conv2_weight_array[0][2][4][2] <= 18'b000000000000111011;\
    conv2_weight_array[0][2][4][3] <= 18'b100000000000010111;\
    conv2_weight_array[0][2][4][4] <= 18'b100000000001110101;\
    conv2_weight_array[0][3][0][0] <= 18'b000000000001111110;\
    conv2_weight_array[0][3][0][1] <= 18'b100000000001101001;\
    conv2_weight_array[0][3][0][2] <= 18'b100000000110000001;\
    conv2_weight_array[0][3][0][3] <= 18'b100000000100110010;\
    conv2_weight_array[0][3][0][4] <= 18'b000000000011001101;\
    conv2_weight_array[0][3][1][0] <= 18'b000000000101001000;\
    conv2_weight_array[0][3][1][1] <= 18'b100000000000001101;\
    conv2_weight_array[0][3][1][2] <= 18'b100000000010100100;\
    conv2_weight_array[0][3][1][3] <= 18'b100000000011000110;\
    conv2_weight_array[0][3][1][4] <= 18'b100000000011010100;\
    conv2_weight_array[0][3][2][0] <= 18'b000000000100101110;\
    conv2_weight_array[0][3][2][1] <= 18'b000000000000000001;\
    conv2_weight_array[0][3][2][2] <= 18'b100000000000011001;\
    conv2_weight_array[0][3][2][3] <= 18'b000000000000010011;\
    conv2_weight_array[0][3][2][4] <= 18'b000000000000000111;\
    conv2_weight_array[0][3][3][0] <= 18'b100000000001000010;\
    conv2_weight_array[0][3][3][1] <= 18'b100000000001110010;\
    conv2_weight_array[0][3][3][2] <= 18'b100000000000110101;\
    conv2_weight_array[0][3][3][3] <= 18'b100000000001110111;\
    conv2_weight_array[0][3][3][4] <= 18'b000000000001100100;\
    conv2_weight_array[0][3][4][0] <= 18'b100000000010010000;\
    conv2_weight_array[0][3][4][1] <= 18'b100000000001000101;\
    conv2_weight_array[0][3][4][2] <= 18'b100000000001001000;\
    conv2_weight_array[0][3][4][3] <= 18'b100000000010110110;\
    conv2_weight_array[0][3][4][4] <= 18'b000000000000011111;\
    conv2_weight_array[0][4][0][0] <= 18'b000000000010111000;\
    conv2_weight_array[0][4][0][1] <= 18'b000000000110100001;\
    conv2_weight_array[0][4][0][2] <= 18'b000000000101010111;\
    conv2_weight_array[0][4][0][3] <= 18'b000000000011011000;\
    conv2_weight_array[0][4][0][4] <= 18'b000000000001111001;\
    conv2_weight_array[0][4][1][0] <= 18'b100000000100000101;\
    conv2_weight_array[0][4][1][1] <= 18'b100000000100100000;\
    conv2_weight_array[0][4][1][2] <= 18'b100000001001110000;\
    conv2_weight_array[0][4][1][3] <= 18'b100000001011110011;\
    conv2_weight_array[0][4][1][4] <= 18'b100000001010110110;\
    conv2_weight_array[0][4][2][0] <= 18'b100000001011000101;\
    conv2_weight_array[0][4][2][1] <= 18'b100000001011110010;\
    conv2_weight_array[0][4][2][2] <= 18'b100000001000111100;\
    conv2_weight_array[0][4][2][3] <= 18'b100000000001110001;\
    conv2_weight_array[0][4][2][4] <= 18'b000000000010011010;\
    conv2_weight_array[0][4][3][0] <= 18'b100000000110001101;\
    conv2_weight_array[0][4][3][1] <= 18'b100000000100111011;\
    conv2_weight_array[0][4][3][2] <= 18'b100000000110110111;\
    conv2_weight_array[0][4][3][3] <= 18'b100000000101100011;\
    conv2_weight_array[0][4][3][4] <= 18'b000000000010000011;\
    conv2_weight_array[0][4][4][0] <= 18'b000000000110111101;\
    conv2_weight_array[0][4][4][1] <= 18'b000000000110101101;\
    conv2_weight_array[0][4][4][2] <= 18'b000000000001111110;\
    conv2_weight_array[0][4][4][3] <= 18'b100000000101111011;\
    conv2_weight_array[0][4][4][4] <= 18'b100000000100100001;\
    conv2_weight_array[0][5][0][0] <= 18'b100000000001111011;\
    conv2_weight_array[0][5][0][1] <= 18'b100000000001100111;\
    conv2_weight_array[0][5][0][2] <= 18'b100000000011011111;\
    conv2_weight_array[0][5][0][3] <= 18'b100000000110010000;\
    conv2_weight_array[0][5][0][4] <= 18'b100000000011100000;\
    conv2_weight_array[0][5][1][0] <= 18'b100000000011110000;\
    conv2_weight_array[0][5][1][1] <= 18'b000000000101111010;\
    conv2_weight_array[0][5][1][2] <= 18'b000000000101011101;\
    conv2_weight_array[0][5][1][3] <= 18'b100000000100111011;\
    conv2_weight_array[0][5][1][4] <= 18'b100000000101110010;\
    conv2_weight_array[0][5][2][0] <= 18'b000000000000010011;\
    conv2_weight_array[0][5][2][1] <= 18'b000000000101000000;\
    conv2_weight_array[0][5][2][2] <= 18'b000000000110111000;\
    conv2_weight_array[0][5][2][3] <= 18'b000000000101001000;\
    conv2_weight_array[0][5][2][4] <= 18'b000000000101010000;\
    conv2_weight_array[0][5][3][0] <= 18'b000000001000011011;\
    conv2_weight_array[0][5][3][1] <= 18'b000000001010010101;\
    conv2_weight_array[0][5][3][2] <= 18'b000000000110011110;\
    conv2_weight_array[0][5][3][3] <= 18'b000000000100100111;\
    conv2_weight_array[0][5][3][4] <= 18'b100000000001101111;\
    conv2_weight_array[0][5][4][0] <= 18'b100000000011010001;\
    conv2_weight_array[0][5][4][1] <= 18'b000000000001011011;\
    conv2_weight_array[0][5][4][2] <= 18'b100000000010010010;\
    conv2_weight_array[0][5][4][3] <= 18'b100000000000101000;\
    conv2_weight_array[0][5][4][4] <= 18'b100000000010010011;\
    conv2_weight_array[1][0][0][0] <= 18'b100000000101000100;\
    conv2_weight_array[1][0][0][1] <= 18'b100000000010001110;\
    conv2_weight_array[1][0][0][2] <= 18'b100000000010001111;\
    conv2_weight_array[1][0][0][3] <= 18'b000000000000000010;\
    conv2_weight_array[1][0][0][4] <= 18'b100000000000000010;\
    conv2_weight_array[1][0][1][0] <= 18'b100000000010101111;\
    conv2_weight_array[1][0][1][1] <= 18'b100000000010010011;\
    conv2_weight_array[1][0][1][2] <= 18'b100000000001100111;\
    conv2_weight_array[1][0][1][3] <= 18'b000000000001010111;\
    conv2_weight_array[1][0][1][4] <= 18'b000000000010100010;\
    conv2_weight_array[1][0][2][0] <= 18'b000000000001101000;\
    conv2_weight_array[1][0][2][1] <= 18'b000000000001010011;\
    conv2_weight_array[1][0][2][2] <= 18'b100000000100100010;\
    conv2_weight_array[1][0][2][3] <= 18'b000000000010001101;\
    conv2_weight_array[1][0][2][4] <= 18'b000000001010111110;\
    conv2_weight_array[1][0][3][0] <= 18'b000000000111100100;\
    conv2_weight_array[1][0][3][1] <= 18'b000000000001011101;\
    conv2_weight_array[1][0][3][2] <= 18'b100000000100000000;\
    conv2_weight_array[1][0][3][3] <= 18'b100000000110101011;\
    conv2_weight_array[1][0][3][4] <= 18'b000000001000000101;\
    conv2_weight_array[1][0][4][0] <= 18'b000000000110011101;\
    conv2_weight_array[1][0][4][1] <= 18'b100000000001001111;\
    conv2_weight_array[1][0][4][2] <= 18'b100000000011111100;\
    conv2_weight_array[1][0][4][3] <= 18'b000000000001000110;\
    conv2_weight_array[1][0][4][4] <= 18'b000000000100110110;\
    conv2_weight_array[1][1][0][0] <= 18'b000000000010001010;\
    conv2_weight_array[1][1][0][1] <= 18'b100000000010100100;\
    conv2_weight_array[1][1][0][2] <= 18'b100000000111010111;\
    conv2_weight_array[1][1][0][3] <= 18'b100000000001100011;\
    conv2_weight_array[1][1][0][4] <= 18'b000000000000000100;\
    conv2_weight_array[1][1][1][0] <= 18'b000000000100010101;\
    conv2_weight_array[1][1][1][1] <= 18'b100000000001001011;\
    conv2_weight_array[1][1][1][2] <= 18'b100000000011001101;\
    conv2_weight_array[1][1][1][3] <= 18'b100000000001010010;\
    conv2_weight_array[1][1][1][4] <= 18'b100000000001000001;\
    conv2_weight_array[1][1][2][0] <= 18'b100000000101110001;\
    conv2_weight_array[1][1][2][1] <= 18'b100000000010010111;\
    conv2_weight_array[1][1][2][2] <= 18'b000000000000010100;\
    conv2_weight_array[1][1][2][3] <= 18'b100000000010101101;\
    conv2_weight_array[1][1][2][4] <= 18'b000000000001111010;\
    conv2_weight_array[1][1][3][0] <= 18'b100000000010011111;\
    conv2_weight_array[1][1][3][1] <= 18'b000000000100101000;\
    conv2_weight_array[1][1][3][2] <= 18'b000000000010000010;\
    conv2_weight_array[1][1][3][3] <= 18'b100000001000110010;\
    conv2_weight_array[1][1][3][4] <= 18'b100000000010000110;\
    conv2_weight_array[1][1][4][0] <= 18'b000000000011010010;\
    conv2_weight_array[1][1][4][1] <= 18'b000000000010000100;\
    conv2_weight_array[1][1][4][2] <= 18'b000000001000000011;\
    conv2_weight_array[1][1][4][3] <= 18'b000000000001110100;\
    conv2_weight_array[1][1][4][4] <= 18'b000000000010101100;\
    conv2_weight_array[1][2][0][0] <= 18'b100000000000111100;\
    conv2_weight_array[1][2][0][1] <= 18'b100000000001110111;\
    conv2_weight_array[1][2][0][2] <= 18'b000000000000101101;\
    conv2_weight_array[1][2][0][3] <= 18'b000000000001000011;\
    conv2_weight_array[1][2][0][4] <= 18'b100000000001001101;\
    conv2_weight_array[1][2][1][0] <= 18'b100000000010011001;\
    conv2_weight_array[1][2][1][1] <= 18'b100000000000010110;\
    conv2_weight_array[1][2][1][2] <= 18'b000000000000010101;\
    conv2_weight_array[1][2][1][3] <= 18'b000000000010011011;\
    conv2_weight_array[1][2][1][4] <= 18'b000000000010001001;\
    conv2_weight_array[1][2][2][0] <= 18'b100000000001000100;\
    conv2_weight_array[1][2][2][1] <= 18'b000000000000000010;\
    conv2_weight_array[1][2][2][2] <= 18'b000000000100010101;\
    conv2_weight_array[1][2][2][3] <= 18'b000000000111011100;\
    conv2_weight_array[1][2][2][4] <= 18'b000000000111101101;\
    conv2_weight_array[1][2][3][0] <= 18'b000000000010011110;\
    conv2_weight_array[1][2][3][1] <= 18'b100000000001111000;\
    conv2_weight_array[1][2][3][2] <= 18'b100000000100010001;\
    conv2_weight_array[1][2][3][3] <= 18'b100000000001101100;\
    conv2_weight_array[1][2][3][4] <= 18'b000000000101010101;\
    conv2_weight_array[1][2][4][0] <= 18'b000000000001001100;\
    conv2_weight_array[1][2][4][1] <= 18'b100000000101110001;\
    conv2_weight_array[1][2][4][2] <= 18'b100000000110001110;\
    conv2_weight_array[1][2][4][3] <= 18'b100000000101101011;\
    conv2_weight_array[1][2][4][4] <= 18'b100000000010000011;\
    conv2_weight_array[1][3][0][0] <= 18'b100000000000010101;\
    conv2_weight_array[1][3][0][1] <= 18'b000000000000100100;\
    conv2_weight_array[1][3][0][2] <= 18'b000000000011011100;\
    conv2_weight_array[1][3][0][3] <= 18'b000000000010101110;\
    conv2_weight_array[1][3][0][4] <= 18'b000000000000100110;\
    conv2_weight_array[1][3][1][0] <= 18'b100000000010011010;\
    conv2_weight_array[1][3][1][1] <= 18'b100000000000110011;\
    conv2_weight_array[1][3][1][2] <= 18'b000000000010110000;\
    conv2_weight_array[1][3][1][3] <= 18'b000000000011011010;\
    conv2_weight_array[1][3][1][4] <= 18'b000000000100100000;\
    conv2_weight_array[1][3][2][0] <= 18'b100000000010000111;\
    conv2_weight_array[1][3][2][1] <= 18'b100000000010010101;\
    conv2_weight_array[1][3][2][2] <= 18'b000000000100000010;\
    conv2_weight_array[1][3][2][3] <= 18'b000000000011110101;\
    conv2_weight_array[1][3][2][4] <= 18'b000000000011000000;\
    conv2_weight_array[1][3][3][0] <= 18'b100000000001001010;\
    conv2_weight_array[1][3][3][1] <= 18'b100000000011111010;\
    conv2_weight_array[1][3][3][2] <= 18'b100000000001101001;\
    conv2_weight_array[1][3][3][3] <= 18'b000000000000001010;\
    conv2_weight_array[1][3][3][4] <= 18'b100000000010001001;\
    conv2_weight_array[1][3][4][0] <= 18'b100000000001100001;\
    conv2_weight_array[1][3][4][1] <= 18'b100000000110000100;\
    conv2_weight_array[1][3][4][2] <= 18'b100000000101010111;\
    conv2_weight_array[1][3][4][3] <= 18'b100000000011101111;\
    conv2_weight_array[1][3][4][4] <= 18'b100000000010101010;\
    conv2_weight_array[1][4][0][0] <= 18'b000000000010011001;\
    conv2_weight_array[1][4][0][1] <= 18'b000000000001001101;\
    conv2_weight_array[1][4][0][2] <= 18'b000000000101100111;\
    conv2_weight_array[1][4][0][3] <= 18'b000000000001010110;\
    conv2_weight_array[1][4][0][4] <= 18'b100000000010111101;\
    conv2_weight_array[1][4][1][0] <= 18'b000000000001000000;\
    conv2_weight_array[1][4][1][1] <= 18'b000000000001010110;\
    conv2_weight_array[1][4][1][2] <= 18'b000000000110101100;\
    conv2_weight_array[1][4][1][3] <= 18'b000000000110001010;\
    conv2_weight_array[1][4][1][4] <= 18'b100000000000100001;\
    conv2_weight_array[1][4][2][0] <= 18'b100000000010001001;\
    conv2_weight_array[1][4][2][1] <= 18'b100000000000111000;\
    conv2_weight_array[1][4][2][2] <= 18'b100000000110101001;\
    conv2_weight_array[1][4][2][3] <= 18'b100000000101010001;\
    conv2_weight_array[1][4][2][4] <= 18'b100000000100010010;\
    conv2_weight_array[1][4][3][0] <= 18'b100000000001011010;\
    conv2_weight_array[1][4][3][1] <= 18'b100000000000000110;\
    conv2_weight_array[1][4][3][2] <= 18'b100000000111111011;\
    conv2_weight_array[1][4][3][3] <= 18'b100000001001000110;\
    conv2_weight_array[1][4][3][4] <= 18'b100000000110100110;\
    conv2_weight_array[1][4][4][0] <= 18'b000000000011000101;\
    conv2_weight_array[1][4][4][1] <= 18'b000000000011100100;\
    conv2_weight_array[1][4][4][2] <= 18'b100000000101111000;\
    conv2_weight_array[1][4][4][3] <= 18'b100000001000001001;\
    conv2_weight_array[1][4][4][4] <= 18'b100000000000001010;\
    conv2_weight_array[1][5][0][0] <= 18'b000000000001111100;\
    conv2_weight_array[1][5][0][1] <= 18'b000000000011010010;\
    conv2_weight_array[1][5][0][2] <= 18'b100000000001001000;\
    conv2_weight_array[1][5][0][3] <= 18'b000000000001100011;\
    conv2_weight_array[1][5][0][4] <= 18'b000000000001011001;\
    conv2_weight_array[1][5][1][0] <= 18'b000000000001001111;\
    conv2_weight_array[1][5][1][1] <= 18'b100000000001101000;\
    conv2_weight_array[1][5][1][2] <= 18'b100000000100001111;\
    conv2_weight_array[1][5][1][3] <= 18'b000000000000011000;\
    conv2_weight_array[1][5][1][4] <= 18'b000000000010001100;\
    conv2_weight_array[1][5][2][0] <= 18'b100000000000010011;\
    conv2_weight_array[1][5][2][1] <= 18'b000000000010010010;\
    conv2_weight_array[1][5][2][2] <= 18'b000000000001000101;\
    conv2_weight_array[1][5][2][3] <= 18'b100000000010100101;\
    conv2_weight_array[1][5][2][4] <= 18'b100000000111010011;\
    conv2_weight_array[1][5][3][0] <= 18'b000000000010000101;\
    conv2_weight_array[1][5][3][1] <= 18'b000000000001111100;\
    conv2_weight_array[1][5][3][2] <= 18'b000000000001011010;\
    conv2_weight_array[1][5][3][3] <= 18'b100000000100101001;\
    conv2_weight_array[1][5][3][4] <= 18'b100000001001001110;\
    conv2_weight_array[1][5][4][0] <= 18'b100000000010000111;\
    conv2_weight_array[1][5][4][1] <= 18'b000000000011001011;\
    conv2_weight_array[1][5][4][2] <= 18'b000000001100000101;\
    conv2_weight_array[1][5][4][3] <= 18'b000000000110011011;\
    conv2_weight_array[1][5][4][4] <= 18'b100000000100000001;\
    conv2_weight_array[2][0][0][0] <= 18'b000000000000101100;\
    conv2_weight_array[2][0][0][1] <= 18'b000000000001110110;\
    conv2_weight_array[2][0][0][2] <= 18'b000000000000000100;\
    conv2_weight_array[2][0][0][3] <= 18'b000000000011010000;\
    conv2_weight_array[2][0][0][4] <= 18'b100000000100011110;\
    conv2_weight_array[2][0][1][0] <= 18'b100000000100010011;\
    conv2_weight_array[2][0][1][1] <= 18'b100000000010111101;\
    conv2_weight_array[2][0][1][2] <= 18'b100000000011111110;\
    conv2_weight_array[2][0][1][3] <= 18'b100000000000001010;\
    conv2_weight_array[2][0][1][4] <= 18'b100000000011011110;\
    conv2_weight_array[2][0][2][0] <= 18'b100000000011100110;\
    conv2_weight_array[2][0][2][1] <= 18'b100000000000010011;\
    conv2_weight_array[2][0][2][2] <= 18'b100000000001001110;\
    conv2_weight_array[2][0][2][3] <= 18'b100000000010010101;\
    conv2_weight_array[2][0][2][4] <= 18'b100000000011000011;\
    conv2_weight_array[2][0][3][0] <= 18'b100000000101111011;\
    conv2_weight_array[2][0][3][1] <= 18'b100000000010010000;\
    conv2_weight_array[2][0][3][2] <= 18'b000000000000101111;\
    conv2_weight_array[2][0][3][3] <= 18'b100000000000001111;\
    conv2_weight_array[2][0][3][4] <= 18'b100000000001000111;\
    conv2_weight_array[2][0][4][0] <= 18'b100000000010100101;\
    conv2_weight_array[2][0][4][1] <= 18'b100000000000010110;\
    conv2_weight_array[2][0][4][2] <= 18'b000000000001111101;\
    conv2_weight_array[2][0][4][3] <= 18'b100000000010010110;\
    conv2_weight_array[2][0][4][4] <= 18'b100000000010111010;\
    conv2_weight_array[2][1][0][0] <= 18'b100000000100011001;\
    conv2_weight_array[2][1][0][1] <= 18'b100000000010100110;\
    conv2_weight_array[2][1][0][2] <= 18'b100000000010000100;\
    conv2_weight_array[2][1][0][3] <= 18'b000000000001010011;\
    conv2_weight_array[2][1][0][4] <= 18'b100000000001000110;\
    conv2_weight_array[2][1][1][0] <= 18'b000000000010000111;\
    conv2_weight_array[2][1][1][1] <= 18'b000000000100110111;\
    conv2_weight_array[2][1][1][2] <= 18'b000000000010110101;\
    conv2_weight_array[2][1][1][3] <= 18'b000000000110011000;\
    conv2_weight_array[2][1][1][4] <= 18'b100000000111000010;\
    conv2_weight_array[2][1][2][0] <= 18'b100000000000101111;\
    conv2_weight_array[2][1][2][1] <= 18'b000000000011011010;\
    conv2_weight_array[2][1][2][2] <= 18'b000000000010000010;\
    conv2_weight_array[2][1][2][3] <= 18'b100000000010101111;\
    conv2_weight_array[2][1][2][4] <= 18'b100000000101011011;\
    conv2_weight_array[2][1][3][0] <= 18'b000000000001001100;\
    conv2_weight_array[2][1][3][1] <= 18'b000000000100100110;\
    conv2_weight_array[2][1][3][2] <= 18'b000000000111000100;\
    conv2_weight_array[2][1][3][3] <= 18'b000000000000100110;\
    conv2_weight_array[2][1][3][4] <= 18'b100000000000110110;\
    conv2_weight_array[2][1][4][0] <= 18'b000000000001011000;\
    conv2_weight_array[2][1][4][1] <= 18'b000000000010000000;\
    conv2_weight_array[2][1][4][2] <= 18'b000000000100010011;\
    conv2_weight_array[2][1][4][3] <= 18'b100000000110011000;\
    conv2_weight_array[2][1][4][4] <= 18'b100000000011100011;\
    conv2_weight_array[2][2][0][0] <= 18'b000000000001100100;\
    conv2_weight_array[2][2][0][1] <= 18'b100000000001101011;\
    conv2_weight_array[2][2][0][2] <= 18'b000000000000110001;\
    conv2_weight_array[2][2][0][3] <= 18'b000000000000110000;\
    conv2_weight_array[2][2][0][4] <= 18'b000000000010001001;\
    conv2_weight_array[2][2][1][0] <= 18'b000000000010101011;\
    conv2_weight_array[2][2][1][1] <= 18'b000000000001000010;\
    conv2_weight_array[2][2][1][2] <= 18'b100000000000010011;\
    conv2_weight_array[2][2][1][3] <= 18'b100000000001100001;\
    conv2_weight_array[2][2][1][4] <= 18'b000000000010110111;\
    conv2_weight_array[2][2][2][0] <= 18'b000000000001100111;\
    conv2_weight_array[2][2][2][1] <= 18'b000000000000101110;\
    conv2_weight_array[2][2][2][2] <= 18'b100000000000101000;\
    conv2_weight_array[2][2][2][3] <= 18'b100000000010111111;\
    conv2_weight_array[2][2][2][4] <= 18'b100000000001000000;\
    conv2_weight_array[2][2][3][0] <= 18'b000000000011000000;\
    conv2_weight_array[2][2][3][1] <= 18'b000000000011100011;\
    conv2_weight_array[2][2][3][2] <= 18'b100000000010000001;\
    conv2_weight_array[2][2][3][3] <= 18'b100000000010100110;\
    conv2_weight_array[2][2][3][4] <= 18'b000000000010010011;\
    conv2_weight_array[2][2][4][0] <= 18'b000000000101110101;\
    conv2_weight_array[2][2][4][1] <= 18'b000000000001100000;\
    conv2_weight_array[2][2][4][2] <= 18'b100000000000100100;\
    conv2_weight_array[2][2][4][3] <= 18'b100000000010100101;\
    conv2_weight_array[2][2][4][4] <= 18'b000000000100101000;\
    conv2_weight_array[2][3][0][0] <= 18'b000000000000110100;\
    conv2_weight_array[2][3][0][1] <= 18'b100000000000111111;\
    conv2_weight_array[2][3][0][2] <= 18'b100000000001100110;\
    conv2_weight_array[2][3][0][3] <= 18'b000000000001101000;\
    conv2_weight_array[2][3][0][4] <= 18'b000000000010100110;\
    conv2_weight_array[2][3][1][0] <= 18'b000000000001111001;\
    conv2_weight_array[2][3][1][1] <= 18'b000000000010011000;\
    conv2_weight_array[2][3][1][2] <= 18'b100000000000000100;\
    conv2_weight_array[2][3][1][3] <= 18'b100000000010111110;\
    conv2_weight_array[2][3][1][4] <= 18'b100000000001010011;\
    conv2_weight_array[2][3][2][0] <= 18'b000000000010100100;\
    conv2_weight_array[2][3][2][1] <= 18'b000000000010100010;\
    conv2_weight_array[2][3][2][2] <= 18'b100000000010000101;\
    conv2_weight_array[2][3][2][3] <= 18'b100000000011001101;\
    conv2_weight_array[2][3][2][4] <= 18'b000000000001111100;\
    conv2_weight_array[2][3][3][0] <= 18'b000000000101110001;\
    conv2_weight_array[2][3][3][1] <= 18'b000000000101001000;\
    conv2_weight_array[2][3][3][2] <= 18'b100000000010111000;\
    conv2_weight_array[2][3][3][3] <= 18'b100000000110111001;\
    conv2_weight_array[2][3][3][4] <= 18'b000000000110010001;\
    conv2_weight_array[2][3][4][0] <= 18'b000000000111011011;\
    conv2_weight_array[2][3][4][1] <= 18'b000000000101101000;\
    conv2_weight_array[2][3][4][2] <= 18'b100000000011000110;\
    conv2_weight_array[2][3][4][3] <= 18'b100000000011001011;\
    conv2_weight_array[2][3][4][4] <= 18'b000000000010100111;\
    conv2_weight_array[2][4][0][0] <= 18'b100000000100101101;\
    conv2_weight_array[2][4][0][1] <= 18'b100000000010110010;\
    conv2_weight_array[2][4][0][2] <= 18'b000000000000100101;\
    conv2_weight_array[2][4][0][3] <= 18'b000000000001110000;\
    conv2_weight_array[2][4][0][4] <= 18'b000000000100101111;\
    conv2_weight_array[2][4][1][0] <= 18'b000000000011101101;\
    conv2_weight_array[2][4][1][1] <= 18'b000000000010000001;\
    conv2_weight_array[2][4][1][2] <= 18'b100000000000010011;\
    conv2_weight_array[2][4][1][3] <= 18'b100000000000011110;\
    conv2_weight_array[2][4][1][4] <= 18'b100000000001100001;\
    conv2_weight_array[2][4][2][0] <= 18'b000000001000011100;\
    conv2_weight_array[2][4][2][1] <= 18'b000000000101000101;\
    conv2_weight_array[2][4][2][2] <= 18'b000000000010000001;\
    conv2_weight_array[2][4][2][3] <= 18'b100000000001001110;\
    conv2_weight_array[2][4][2][4] <= 18'b100000000111111100;\
    conv2_weight_array[2][4][3][0] <= 18'b000000000101000111;\
    conv2_weight_array[2][4][3][1] <= 18'b000000000001000110;\
    conv2_weight_array[2][4][3][2] <= 18'b000000000001101100;\
    conv2_weight_array[2][4][3][3] <= 18'b000000000000001101;\
    conv2_weight_array[2][4][3][4] <= 18'b100000000011011010;\
    conv2_weight_array[2][4][4][0] <= 18'b000000000110111001;\
    conv2_weight_array[2][4][4][1] <= 18'b000000000000000000;\
    conv2_weight_array[2][4][4][2] <= 18'b000000000010001101;\
    conv2_weight_array[2][4][4][3] <= 18'b000000000000110101;\
    conv2_weight_array[2][4][4][4] <= 18'b100000000000000110;\
    conv2_weight_array[2][5][0][0] <= 18'b100000000100101110;\
    conv2_weight_array[2][5][0][1] <= 18'b000000000001010100;\
    conv2_weight_array[2][5][0][2] <= 18'b100000000000101101;\
    conv2_weight_array[2][5][0][3] <= 18'b000000000010001000;\
    conv2_weight_array[2][5][0][4] <= 18'b000000000000110000;\
    conv2_weight_array[2][5][1][0] <= 18'b000000000000000000;\
    conv2_weight_array[2][5][1][1] <= 18'b100000000000111011;\
    conv2_weight_array[2][5][1][2] <= 18'b100000000000011001;\
    conv2_weight_array[2][5][1][3] <= 18'b000000000010101000;\
    conv2_weight_array[2][5][1][4] <= 18'b000000000000010001;\
    conv2_weight_array[2][5][2][0] <= 18'b100000000010100101;\
    conv2_weight_array[2][5][2][1] <= 18'b000000000011010000;\
    conv2_weight_array[2][5][2][2] <= 18'b100000000010100111;\
    conv2_weight_array[2][5][2][3] <= 18'b100000000001010101;\
    conv2_weight_array[2][5][2][4] <= 18'b100000000001001111;\
    conv2_weight_array[2][5][3][0] <= 18'b100000000001001001;\
    conv2_weight_array[2][5][3][1] <= 18'b100000000001011100;\
    conv2_weight_array[2][5][3][2] <= 18'b100000000011000000;\
    conv2_weight_array[2][5][3][3] <= 18'b000000000000100001;\
    conv2_weight_array[2][5][3][4] <= 18'b100000000001111010;\
    conv2_weight_array[2][5][4][0] <= 18'b100000000000010111;\
    conv2_weight_array[2][5][4][1] <= 18'b100000000010010100;\
    conv2_weight_array[2][5][4][2] <= 18'b000000000100001101;\
    conv2_weight_array[2][5][4][3] <= 18'b000000000010100110;\
    conv2_weight_array[2][5][4][4] <= 18'b100000000101101100;\
    conv2_weight_array[3][0][0][0] <= 18'b000000000001000110;\
    conv2_weight_array[3][0][0][1] <= 18'b000000000000010110;\
    conv2_weight_array[3][0][0][2] <= 18'b000000000000100100;\
    conv2_weight_array[3][0][0][3] <= 18'b000000000011000000;\
    conv2_weight_array[3][0][0][4] <= 18'b000000000011111000;\
    conv2_weight_array[3][0][1][0] <= 18'b000000000000011011;\
    conv2_weight_array[3][0][1][1] <= 18'b100000000010000010;\
    conv2_weight_array[3][0][1][2] <= 18'b100000000101010111;\
    conv2_weight_array[3][0][1][3] <= 18'b100000000010110110;\
    conv2_weight_array[3][0][1][4] <= 18'b000000000010100001;\
    conv2_weight_array[3][0][2][0] <= 18'b000000000000110000;\
    conv2_weight_array[3][0][2][1] <= 18'b100000000000001110;\
    conv2_weight_array[3][0][2][2] <= 18'b100000000100101100;\
    conv2_weight_array[3][0][2][3] <= 18'b100000000010100100;\
    conv2_weight_array[3][0][2][4] <= 18'b100000000000001111;\
    conv2_weight_array[3][0][3][0] <= 18'b000000000010000100;\
    conv2_weight_array[3][0][3][1] <= 18'b100000000010100010;\
    conv2_weight_array[3][0][3][2] <= 18'b100000000111010011;\
    conv2_weight_array[3][0][3][3] <= 18'b100000000101110001;\
    conv2_weight_array[3][0][3][4] <= 18'b000000000010001101;\
    conv2_weight_array[3][0][4][0] <= 18'b100000000011110010;\
    conv2_weight_array[3][0][4][1] <= 18'b100000000101011111;\
    conv2_weight_array[3][0][4][2] <= 18'b100000001001011001;\
    conv2_weight_array[3][0][4][3] <= 18'b000000000001000010;\
    conv2_weight_array[3][0][4][4] <= 18'b000000000100001010;\
    conv2_weight_array[3][1][0][0] <= 18'b000000000011100101;\
    conv2_weight_array[3][1][0][1] <= 18'b100000000010010110;\
    conv2_weight_array[3][1][0][2] <= 18'b100000000000011011;\
    conv2_weight_array[3][1][0][3] <= 18'b000000000011111001;\
    conv2_weight_array[3][1][0][4] <= 18'b000000000001001101;\
    conv2_weight_array[3][1][1][0] <= 18'b000000000001010111;\
    conv2_weight_array[3][1][1][1] <= 18'b100000000101010101;\
    conv2_weight_array[3][1][1][2] <= 18'b100000000011111111;\
    conv2_weight_array[3][1][1][3] <= 18'b000000000011110101;\
    conv2_weight_array[3][1][1][4] <= 18'b000000000100100001;\
    conv2_weight_array[3][1][2][0] <= 18'b100000000010011001;\
    conv2_weight_array[3][1][2][1] <= 18'b100000000010111010;\
    conv2_weight_array[3][1][2][2] <= 18'b100000000000111110;\
    conv2_weight_array[3][1][2][3] <= 18'b000000000100110011;\
    conv2_weight_array[3][1][2][4] <= 18'b000000000101000000;\
    conv2_weight_array[3][1][3][0] <= 18'b000000000010011000;\
    conv2_weight_array[3][1][3][1] <= 18'b100000000000010110;\
    conv2_weight_array[3][1][3][2] <= 18'b000000000011111100;\
    conv2_weight_array[3][1][3][3] <= 18'b000000000000001001;\
    conv2_weight_array[3][1][3][4] <= 18'b000000000100000010;\
    conv2_weight_array[3][1][4][0] <= 18'b000000000000100101;\
    conv2_weight_array[3][1][4][1] <= 18'b000000000010110001;\
    conv2_weight_array[3][1][4][2] <= 18'b000000000000100011;\
    conv2_weight_array[3][1][4][3] <= 18'b000000000100001010;\
    conv2_weight_array[3][1][4][4] <= 18'b100000000011001100;\
    conv2_weight_array[3][2][0][0] <= 18'b000000000000011000;\
    conv2_weight_array[3][2][0][1] <= 18'b100000000010101001;\
    conv2_weight_array[3][2][0][2] <= 18'b100000000000110100;\
    conv2_weight_array[3][2][0][3] <= 18'b100000000000011100;\
    conv2_weight_array[3][2][0][4] <= 18'b100000000000011010;\
    conv2_weight_array[3][2][1][0] <= 18'b000000000001110100;\
    conv2_weight_array[3][2][1][1] <= 18'b100000000001000101;\
    conv2_weight_array[3][2][1][2] <= 18'b000000000000101100;\
    conv2_weight_array[3][2][1][3] <= 18'b000000000000011010;\
    conv2_weight_array[3][2][1][4] <= 18'b000000000001110110;\
    conv2_weight_array[3][2][2][0] <= 18'b000000000000111001;\
    conv2_weight_array[3][2][2][1] <= 18'b100000000100001101;\
    conv2_weight_array[3][2][2][2] <= 18'b000000000010101010;\
    conv2_weight_array[3][2][2][3] <= 18'b000000000100001111;\
    conv2_weight_array[3][2][2][4] <= 18'b100000000001010101;\
    conv2_weight_array[3][2][3][0] <= 18'b100000000000000010;\
    conv2_weight_array[3][2][3][1] <= 18'b100000000010000011;\
    conv2_weight_array[3][2][3][2] <= 18'b000000000000100101;\
    conv2_weight_array[3][2][3][3] <= 18'b000000000100001011;\
    conv2_weight_array[3][2][3][4] <= 18'b000000000000011111;\
    conv2_weight_array[3][2][4][0] <= 18'b100000000010101110;\
    conv2_weight_array[3][2][4][1] <= 18'b000000000000110111;\
    conv2_weight_array[3][2][4][2] <= 18'b000000000100110100;\
    conv2_weight_array[3][2][4][3] <= 18'b000000000100111010;\
    conv2_weight_array[3][2][4][4] <= 18'b100000000000000110;\
    conv2_weight_array[3][3][0][0] <= 18'b000000000000011001;\
    conv2_weight_array[3][3][0][1] <= 18'b100000000000001110;\
    conv2_weight_array[3][3][0][2] <= 18'b100000000100011000;\
    conv2_weight_array[3][3][0][3] <= 18'b100000000000100000;\
    conv2_weight_array[3][3][0][4] <= 18'b100000000010011100;\
    conv2_weight_array[3][3][1][0] <= 18'b000000000011001001;\
    conv2_weight_array[3][3][1][1] <= 18'b100000000000110100;\
    conv2_weight_array[3][3][1][2] <= 18'b100000000001001101;\
    conv2_weight_array[3][3][1][3] <= 18'b000000000000100111;\
    conv2_weight_array[3][3][1][4] <= 18'b100000000001001010;\
    conv2_weight_array[3][3][2][0] <= 18'b100000000010100111;\
    conv2_weight_array[3][3][2][1] <= 18'b100000000000101100;\
    conv2_weight_array[3][3][2][2] <= 18'b000000000001011101;\
    conv2_weight_array[3][3][2][3] <= 18'b000000000110000101;\
    conv2_weight_array[3][3][2][4] <= 18'b000000000001110000;\
    conv2_weight_array[3][3][3][0] <= 18'b100000000000010111;\
    conv2_weight_array[3][3][3][1] <= 18'b000000000000011100;\
    conv2_weight_array[3][3][3][2] <= 18'b000000000100001000;\
    conv2_weight_array[3][3][3][3] <= 18'b000000000101100000;\
    conv2_weight_array[3][3][3][4] <= 18'b100000000010111011;\
    conv2_weight_array[3][3][4][0] <= 18'b100000000000100101;\
    conv2_weight_array[3][3][4][1] <= 18'b000000000101111011;\
    conv2_weight_array[3][3][4][2] <= 18'b000000000111110100;\
    conv2_weight_array[3][3][4][3] <= 18'b000000000010011110;\
    conv2_weight_array[3][3][4][4] <= 18'b100000000101101010;\
    conv2_weight_array[3][4][0][0] <= 18'b000000000111110000;\
    conv2_weight_array[3][4][0][1] <= 18'b000000000100010010;\
    conv2_weight_array[3][4][0][2] <= 18'b000000000101011010;\
    conv2_weight_array[3][4][0][3] <= 18'b000000000100001100;\
    conv2_weight_array[3][4][0][4] <= 18'b100000000000101001;\
    conv2_weight_array[3][4][1][0] <= 18'b000000000000101111;\
    conv2_weight_array[3][4][1][1] <= 18'b000000000001001010;\
    conv2_weight_array[3][4][1][2] <= 18'b000000000010111100;\
    conv2_weight_array[3][4][1][3] <= 18'b000000000100000110;\
    conv2_weight_array[3][4][1][4] <= 18'b100000001000010010;\
    conv2_weight_array[3][4][2][0] <= 18'b100000000011111101;\
    conv2_weight_array[3][4][2][1] <= 18'b100000000010111001;\
    conv2_weight_array[3][4][2][2] <= 18'b100000000011001101;\
    conv2_weight_array[3][4][2][3] <= 18'b100000000101101001;\
    conv2_weight_array[3][4][2][4] <= 18'b100000000111111111;\
    conv2_weight_array[3][4][3][0] <= 18'b100000010010110111;\
    conv2_weight_array[3][4][3][1] <= 18'b100000000010101001;\
    conv2_weight_array[3][4][3][2] <= 18'b100000000101010111;\
    conv2_weight_array[3][4][3][3] <= 18'b100000000010000100;\
    conv2_weight_array[3][4][3][4] <= 18'b100000000101100000;\
    conv2_weight_array[3][4][4][0] <= 18'b100000001010000001;\
    conv2_weight_array[3][4][4][1] <= 18'b000000000100111000;\
    conv2_weight_array[3][4][4][2] <= 18'b000000000011101001;\
    conv2_weight_array[3][4][4][3] <= 18'b100000000011001111;\
    conv2_weight_array[3][4][4][4] <= 18'b100000000011111101;\
    conv2_weight_array[3][5][0][0] <= 18'b000000000011110110;\
    conv2_weight_array[3][5][0][1] <= 18'b000000000000100111;\
    conv2_weight_array[3][5][0][2] <= 18'b000000000000110101;\
    conv2_weight_array[3][5][0][3] <= 18'b000000000001001010;\
    conv2_weight_array[3][5][0][4] <= 18'b000000000010000011;\
    conv2_weight_array[3][5][1][0] <= 18'b000000000010100000;\
    conv2_weight_array[3][5][1][1] <= 18'b100000000011100101;\
    conv2_weight_array[3][5][1][2] <= 18'b000000000001001100;\
    conv2_weight_array[3][5][1][3] <= 18'b000000000011000101;\
    conv2_weight_array[3][5][1][4] <= 18'b000000001011011101;\
    conv2_weight_array[3][5][2][0] <= 18'b100000000101100110;\
    conv2_weight_array[3][5][2][1] <= 18'b000000000001100010;\
    conv2_weight_array[3][5][2][2] <= 18'b000000000101010000;\
    conv2_weight_array[3][5][2][3] <= 18'b000000001001000111;\
    conv2_weight_array[3][5][2][4] <= 18'b000000000110000111;\
    conv2_weight_array[3][5][3][0] <= 18'b000000000001100001;\
    conv2_weight_array[3][5][3][1] <= 18'b000000000100110101;\
    conv2_weight_array[3][5][3][2] <= 18'b000000000001111011;\
    conv2_weight_array[3][5][3][3] <= 18'b100000000000000001;\
    conv2_weight_array[3][5][3][4] <= 18'b000000000001010000;\
    conv2_weight_array[3][5][4][0] <= 18'b000000000100111100;\
    conv2_weight_array[3][5][4][1] <= 18'b100000000000100000;\
    conv2_weight_array[3][5][4][2] <= 18'b100000000011001001;\
    conv2_weight_array[3][5][4][3] <= 18'b100000000111100000;\
    conv2_weight_array[3][5][4][4] <= 18'b100000000000110010;\
    conv2_weight_array[4][0][0][0] <= 18'b000000000100000110;\
    conv2_weight_array[4][0][0][1] <= 18'b000000000011000111;\
    conv2_weight_array[4][0][0][2] <= 18'b100000000001111000;\
    conv2_weight_array[4][0][0][3] <= 18'b100000000010011100;\
    conv2_weight_array[4][0][0][4] <= 18'b000000000000101100;\
    conv2_weight_array[4][0][1][0] <= 18'b000000000010111000;\
    conv2_weight_array[4][0][1][1] <= 18'b000000000011001010;\
    conv2_weight_array[4][0][1][2] <= 18'b100000000010101100;\
    conv2_weight_array[4][0][1][3] <= 18'b100000000010101111;\
    conv2_weight_array[4][0][1][4] <= 18'b100000000000010110;\
    conv2_weight_array[4][0][2][0] <= 18'b100000000000000010;\
    conv2_weight_array[4][0][2][1] <= 18'b100000000000010010;\
    conv2_weight_array[4][0][2][2] <= 18'b000000000100110010;\
    conv2_weight_array[4][0][2][3] <= 18'b000000000110101010;\
    conv2_weight_array[4][0][2][4] <= 18'b100000000011010110;\
    conv2_weight_array[4][0][3][0] <= 18'b100000001011100100;\
    conv2_weight_array[4][0][3][1] <= 18'b100000000111110110;\
    conv2_weight_array[4][0][3][2] <= 18'b000000000010100101;\
    conv2_weight_array[4][0][3][3] <= 18'b000000001011010001;\
    conv2_weight_array[4][0][3][4] <= 18'b000000000101101111;\
    conv2_weight_array[4][0][4][0] <= 18'b000000000000101011;\
    conv2_weight_array[4][0][4][1] <= 18'b000000000010011010;\
    conv2_weight_array[4][0][4][2] <= 18'b100000000110100001;\
    conv2_weight_array[4][0][4][3] <= 18'b000000000010001000;\
    conv2_weight_array[4][0][4][4] <= 18'b000000000010111001;\
    conv2_weight_array[4][1][0][0] <= 18'b100000000010111001;\
    conv2_weight_array[4][1][0][1] <= 18'b000000000010110110;\
    conv2_weight_array[4][1][0][2] <= 18'b000000000110011111;\
    conv2_weight_array[4][1][0][3] <= 18'b000000000011000111;\
    conv2_weight_array[4][1][0][4] <= 18'b000000000011010000;\
    conv2_weight_array[4][1][1][0] <= 18'b100000000001011000;\
    conv2_weight_array[4][1][1][1] <= 18'b100000000011100100;\
    conv2_weight_array[4][1][1][2] <= 18'b000000000101101111;\
    conv2_weight_array[4][1][1][3] <= 18'b000000000111011110;\
    conv2_weight_array[4][1][1][4] <= 18'b000000000000001010;\
    conv2_weight_array[4][1][2][0] <= 18'b000000000000110110;\
    conv2_weight_array[4][1][2][1] <= 18'b100000000010101110;\
    conv2_weight_array[4][1][2][2] <= 18'b100000000010010010;\
    conv2_weight_array[4][1][2][3] <= 18'b000000000100111100;\
    conv2_weight_array[4][1][2][4] <= 18'b000000000001010000;\
    conv2_weight_array[4][1][3][0] <= 18'b100000000000111110;\
    conv2_weight_array[4][1][3][1] <= 18'b000000000000000101;\
    conv2_weight_array[4][1][3][2] <= 18'b100000000110100111;\
    conv2_weight_array[4][1][3][3] <= 18'b000000000000111111;\
    conv2_weight_array[4][1][3][4] <= 18'b000000000001001110;\
    conv2_weight_array[4][1][4][0] <= 18'b100000000000000011;\
    conv2_weight_array[4][1][4][1] <= 18'b100000000001011110;\
    conv2_weight_array[4][1][4][2] <= 18'b100000000111000111;\
    conv2_weight_array[4][1][4][3] <= 18'b100000000011101010;\
    conv2_weight_array[4][1][4][4] <= 18'b100000000000000110;\
    conv2_weight_array[4][2][0][0] <= 18'b000000000100001101;\
    conv2_weight_array[4][2][0][1] <= 18'b100000000001011110;\
    conv2_weight_array[4][2][0][2] <= 18'b100000000101011000;\
    conv2_weight_array[4][2][0][3] <= 18'b100000000001100110;\
    conv2_weight_array[4][2][0][4] <= 18'b100000000010000100;\
    conv2_weight_array[4][2][1][0] <= 18'b000000000011100101;\
    conv2_weight_array[4][2][1][1] <= 18'b000000000010000110;\
    conv2_weight_array[4][2][1][2] <= 18'b100000000000001001;\
    conv2_weight_array[4][2][1][3] <= 18'b100000000001100111;\
    conv2_weight_array[4][2][1][4] <= 18'b100000000011011111;\
    conv2_weight_array[4][2][2][0] <= 18'b000000000000010001;\
    conv2_weight_array[4][2][2][1] <= 18'b000000000100010101;\
    conv2_weight_array[4][2][2][2] <= 18'b000000000010011100;\
    conv2_weight_array[4][2][2][3] <= 18'b000000000010010001;\
    conv2_weight_array[4][2][2][4] <= 18'b100000000011111001;\
    conv2_weight_array[4][2][3][0] <= 18'b100000000101010111;\
    conv2_weight_array[4][2][3][1] <= 18'b100000000001010001;\
    conv2_weight_array[4][2][3][2] <= 18'b000000000101000001;\
    conv2_weight_array[4][2][3][3] <= 18'b000000001000000110;\
    conv2_weight_array[4][2][3][4] <= 18'b000000000000110011;\
    conv2_weight_array[4][2][4][0] <= 18'b100000000101010000;\
    conv2_weight_array[4][2][4][1] <= 18'b100000000101100110;\
    conv2_weight_array[4][2][4][2] <= 18'b100000000011110110;\
    conv2_weight_array[4][2][4][3] <= 18'b000000000011101001;\
    conv2_weight_array[4][2][4][4] <= 18'b000000000010111111;\
    conv2_weight_array[4][3][0][0] <= 18'b000000000010001001;\
    conv2_weight_array[4][3][0][1] <= 18'b000000000000001111;\
    conv2_weight_array[4][3][0][2] <= 18'b100000000001010111;\
    conv2_weight_array[4][3][0][3] <= 18'b000000000000000011;\
    conv2_weight_array[4][3][0][4] <= 18'b100000000010001100;\
    conv2_weight_array[4][3][1][0] <= 18'b000000000010100101;\
    conv2_weight_array[4][3][1][1] <= 18'b000000000001111110;\
    conv2_weight_array[4][3][1][2] <= 18'b000000000011000100;\
    conv2_weight_array[4][3][1][3] <= 18'b000000000000111110;\
    conv2_weight_array[4][3][1][4] <= 18'b100000000100011100;\
    conv2_weight_array[4][3][2][0] <= 18'b000000000001110000;\
    conv2_weight_array[4][3][2][1] <= 18'b000000000001100000;\
    conv2_weight_array[4][3][2][2] <= 18'b000000000101010010;\
    conv2_weight_array[4][3][2][3] <= 18'b000000000001011110;\
    conv2_weight_array[4][3][2][4] <= 18'b100000000100001101;\
    conv2_weight_array[4][3][3][0] <= 18'b100000000001011100;\
    conv2_weight_array[4][3][3][1] <= 18'b100000000001010000;\
    conv2_weight_array[4][3][3][2] <= 18'b000000000010110011;\
    conv2_weight_array[4][3][3][3] <= 18'b000000000001100110;\
    conv2_weight_array[4][3][3][4] <= 18'b100000000001010101;\
    conv2_weight_array[4][3][4][0] <= 18'b100000000001111110;\
    conv2_weight_array[4][3][4][1] <= 18'b100000000101001100;\
    conv2_weight_array[4][3][4][2] <= 18'b100000000100011011;\
    conv2_weight_array[4][3][4][3] <= 18'b100000000011011010;\
    conv2_weight_array[4][3][4][4] <= 18'b100000000100010111;\
    conv2_weight_array[4][4][0][0] <= 18'b000000000100000110;\
    conv2_weight_array[4][4][0][1] <= 18'b000000000001100101;\
    conv2_weight_array[4][4][0][2] <= 18'b100000000011011110;\
    conv2_weight_array[4][4][0][3] <= 18'b100000000110011111;\
    conv2_weight_array[4][4][0][4] <= 18'b100000000011101101;\
    conv2_weight_array[4][4][1][0] <= 18'b100000001100000101;\
    conv2_weight_array[4][4][1][1] <= 18'b100000000001010110;\
    conv2_weight_array[4][4][1][2] <= 18'b000000000010110010;\
    conv2_weight_array[4][4][1][3] <= 18'b100000000101101101;\
    conv2_weight_array[4][4][1][4] <= 18'b100000000100111100;\
    conv2_weight_array[4][4][2][0] <= 18'b100000000111110111;\
    conv2_weight_array[4][4][2][1] <= 18'b100000000101001010;\
    conv2_weight_array[4][4][2][2] <= 18'b100000000110111001;\
    conv2_weight_array[4][4][2][3] <= 18'b100000000010010111;\
    conv2_weight_array[4][4][2][4] <= 18'b000000000000100001;\
    conv2_weight_array[4][4][3][0] <= 18'b000000000001110111;\
    conv2_weight_array[4][4][3][1] <= 18'b100000000001010001;\
    conv2_weight_array[4][4][3][2] <= 18'b100000001110000010;\
    conv2_weight_array[4][4][3][3] <= 18'b100000001100001000;\
    conv2_weight_array[4][4][3][4] <= 18'b100000000011100010;\
    conv2_weight_array[4][4][4][0] <= 18'b100000000001111000;\
    conv2_weight_array[4][4][4][1] <= 18'b100000000010101110;\
    conv2_weight_array[4][4][4][2] <= 18'b100000001101011101;\
    conv2_weight_array[4][4][4][3] <= 18'b100000000101110111;\
    conv2_weight_array[4][4][4][4] <= 18'b000000000001101010;\
    conv2_weight_array[4][5][0][0] <= 18'b000000000001010100;\
    conv2_weight_array[4][5][0][1] <= 18'b000000000010111100;\
    conv2_weight_array[4][5][0][2] <= 18'b000000000101101111;\
    conv2_weight_array[4][5][0][3] <= 18'b000000001000000011;\
    conv2_weight_array[4][5][0][4] <= 18'b000000000100111101;\
    conv2_weight_array[4][5][1][0] <= 18'b000000000000000001;\
    conv2_weight_array[4][5][1][1] <= 18'b000000000110101101;\
    conv2_weight_array[4][5][1][2] <= 18'b000000000110111000;\
    conv2_weight_array[4][5][1][3] <= 18'b000000001001110001;\
    conv2_weight_array[4][5][1][4] <= 18'b000000000101111100;\
    conv2_weight_array[4][5][2][0] <= 18'b100000000001001100;\
    conv2_weight_array[4][5][2][1] <= 18'b100000000100001111;\
    conv2_weight_array[4][5][2][2] <= 18'b100000000010110110;\
    conv2_weight_array[4][5][2][3] <= 18'b000000000111010100;\
    conv2_weight_array[4][5][2][4] <= 18'b000000000001111100;\
    conv2_weight_array[4][5][3][0] <= 18'b100000000001000010;\
    conv2_weight_array[4][5][3][1] <= 18'b100000000011111000;\
    conv2_weight_array[4][5][3][2] <= 18'b100000000001100011;\
    conv2_weight_array[4][5][3][3] <= 18'b100000000011010100;\
    conv2_weight_array[4][5][3][4] <= 18'b000000000001011000;\
    conv2_weight_array[4][5][4][0] <= 18'b100000000110011101;\
    conv2_weight_array[4][5][4][1] <= 18'b100000000001011100;\
    conv2_weight_array[4][5][4][2] <= 18'b100000000011001010;\
    conv2_weight_array[4][5][4][3] <= 18'b000000000001111000;\
    conv2_weight_array[4][5][4][4] <= 18'b100000000000100101;\
    conv2_weight_array[5][0][0][0] <= 18'b000000000000000101;\
    conv2_weight_array[5][0][0][1] <= 18'b000000000010001011;\
    conv2_weight_array[5][0][0][2] <= 18'b000000000000010000;\
    conv2_weight_array[5][0][0][3] <= 18'b100000000000100110;\
    conv2_weight_array[5][0][0][4] <= 18'b000000000000110001;\
    conv2_weight_array[5][0][1][0] <= 18'b000000000010101001;\
    conv2_weight_array[5][0][1][1] <= 18'b000000000000000011;\
    conv2_weight_array[5][0][1][2] <= 18'b100000000010101100;\
    conv2_weight_array[5][0][1][3] <= 18'b000000000000010000;\
    conv2_weight_array[5][0][1][4] <= 18'b000000000001101100;\
    conv2_weight_array[5][0][2][0] <= 18'b000000000110001010;\
    conv2_weight_array[5][0][2][1] <= 18'b000000000101000000;\
    conv2_weight_array[5][0][2][2] <= 18'b000000000011110110;\
    conv2_weight_array[5][0][2][3] <= 18'b000000000100111100;\
    conv2_weight_array[5][0][2][4] <= 18'b000000000011000110;\
    conv2_weight_array[5][0][3][0] <= 18'b100000000010110011;\
    conv2_weight_array[5][0][3][1] <= 18'b100000000100010101;\
    conv2_weight_array[5][0][3][2] <= 18'b100000000001001011;\
    conv2_weight_array[5][0][3][3] <= 18'b100000000010011110;\
    conv2_weight_array[5][0][3][4] <= 18'b100000000111111010;\
    conv2_weight_array[5][0][4][0] <= 18'b000000000010110110;\
    conv2_weight_array[5][0][4][1] <= 18'b000000000101101001;\
    conv2_weight_array[5][0][4][2] <= 18'b000000000010100001;\
    conv2_weight_array[5][0][4][3] <= 18'b000000000001101111;\
    conv2_weight_array[5][0][4][4] <= 18'b000000000000011001;\
    conv2_weight_array[5][1][0][0] <= 18'b100000000101101100;\
    conv2_weight_array[5][1][0][1] <= 18'b000000000000101111;\
    conv2_weight_array[5][1][0][2] <= 18'b000000000000001110;\
    conv2_weight_array[5][1][0][3] <= 18'b100000000011111101;\
    conv2_weight_array[5][1][0][4] <= 18'b100000000101011101;\
    conv2_weight_array[5][1][1][0] <= 18'b100000000011001101;\
    conv2_weight_array[5][1][1][1] <= 18'b000000000011111101;\
    conv2_weight_array[5][1][1][2] <= 18'b000000000011000101;\
    conv2_weight_array[5][1][1][3] <= 18'b000000000000110110;\
    conv2_weight_array[5][1][1][4] <= 18'b000000000101001001;\
    conv2_weight_array[5][1][2][0] <= 18'b100000000000100111;\
    conv2_weight_array[5][1][2][1] <= 18'b000000000000010100;\
    conv2_weight_array[5][1][2][2] <= 18'b000000000000001000;\
    conv2_weight_array[5][1][2][3] <= 18'b000000000101101010;\
    conv2_weight_array[5][1][2][4] <= 18'b000000001001111001;\
    conv2_weight_array[5][1][3][0] <= 18'b000000000011001000;\
    conv2_weight_array[5][1][3][1] <= 18'b000000000100111111;\
    conv2_weight_array[5][1][3][2] <= 18'b000000000011101101;\
    conv2_weight_array[5][1][3][3] <= 18'b000000000110110011;\
    conv2_weight_array[5][1][3][4] <= 18'b000000000100001111;\
    conv2_weight_array[5][1][4][0] <= 18'b100000000010110100;\
    conv2_weight_array[5][1][4][1] <= 18'b100000001000011110;\
    conv2_weight_array[5][1][4][2] <= 18'b100000000011001111;\
    conv2_weight_array[5][1][4][3] <= 18'b100000000101111110;\
    conv2_weight_array[5][1][4][4] <= 18'b100000000000011110;\
    conv2_weight_array[5][2][0][0] <= 18'b100000000001110110;\
    conv2_weight_array[5][2][0][1] <= 18'b000000000000100111;\
    conv2_weight_array[5][2][0][2] <= 18'b000000000001011000;\
    conv2_weight_array[5][2][0][3] <= 18'b100000000001010011;\
    conv2_weight_array[5][2][0][4] <= 18'b100000000000110001;\
    conv2_weight_array[5][2][1][0] <= 18'b100000000010100110;\
    conv2_weight_array[5][2][1][1] <= 18'b100000000001000111;\
    conv2_weight_array[5][2][1][2] <= 18'b100000000000001110;\
    conv2_weight_array[5][2][1][3] <= 18'b000000000001011000;\
    conv2_weight_array[5][2][1][4] <= 18'b000000000001010001;\
    conv2_weight_array[5][2][2][0] <= 18'b000000000101101010;\
    conv2_weight_array[5][2][2][1] <= 18'b000000000100101010;\
    conv2_weight_array[5][2][2][2] <= 18'b000000000111001001;\
    conv2_weight_array[5][2][2][3] <= 18'b000000000101100101;\
    conv2_weight_array[5][2][2][4] <= 18'b000000000011000001;\
    conv2_weight_array[5][2][3][0] <= 18'b100000000000101110;\
    conv2_weight_array[5][2][3][1] <= 18'b000000000000001110;\
    conv2_weight_array[5][2][3][2] <= 18'b100000000000011110;\
    conv2_weight_array[5][2][3][3] <= 18'b100000000010011000;\
    conv2_weight_array[5][2][3][4] <= 18'b100000000110110110;\
    conv2_weight_array[5][2][4][0] <= 18'b100000000010000110;\
    conv2_weight_array[5][2][4][1] <= 18'b100000000101101010;\
    conv2_weight_array[5][2][4][2] <= 18'b100000000110111110;\
    conv2_weight_array[5][2][4][3] <= 18'b100000001000110111;\
    conv2_weight_array[5][2][4][4] <= 18'b100000000111000110;\
    conv2_weight_array[5][3][0][0] <= 18'b100000000100110111;\
    conv2_weight_array[5][3][0][1] <= 18'b100000000010110000;\
    conv2_weight_array[5][3][0][2] <= 18'b100000000000111000;\
    conv2_weight_array[5][3][0][3] <= 18'b100000000010010000;\
    conv2_weight_array[5][3][0][4] <= 18'b100000000000001000;\
    conv2_weight_array[5][3][1][0] <= 18'b100000000100100011;\
    conv2_weight_array[5][3][1][1] <= 18'b000000000000000010;\
    conv2_weight_array[5][3][1][2] <= 18'b000000000000110101;\
    conv2_weight_array[5][3][1][3] <= 18'b000000000001011110;\
    conv2_weight_array[5][3][1][4] <= 18'b000000000011101101;\
    conv2_weight_array[5][3][2][0] <= 18'b000000000001001000;\
    conv2_weight_array[5][3][2][1] <= 18'b000000000100100000;\
    conv2_weight_array[5][3][2][2] <= 18'b000000000100101011;\
    conv2_weight_array[5][3][2][3] <= 18'b000000000111000110;\
    conv2_weight_array[5][3][2][4] <= 18'b000000000010010011;\
    conv2_weight_array[5][3][3][0] <= 18'b000000000001001011;\
    conv2_weight_array[5][3][3][1] <= 18'b100000000000000101;\
    conv2_weight_array[5][3][3][2] <= 18'b100000000011010111;\
    conv2_weight_array[5][3][3][3] <= 18'b100000000100100010;\
    conv2_weight_array[5][3][3][4] <= 18'b100000000110000011;\
    conv2_weight_array[5][3][4][0] <= 18'b000000000000001111;\
    conv2_weight_array[5][3][4][1] <= 18'b100000000110001100;\
    conv2_weight_array[5][3][4][2] <= 18'b100000000111110100;\
    conv2_weight_array[5][3][4][3] <= 18'b100000000101010100;\
    conv2_weight_array[5][3][4][4] <= 18'b100000000001111001;\
    conv2_weight_array[5][4][0][0] <= 18'b000000000100010110;\
    conv2_weight_array[5][4][0][1] <= 18'b000000000000111111;\
    conv2_weight_array[5][4][0][2] <= 18'b000000000010111010;\
    conv2_weight_array[5][4][0][3] <= 18'b100000000000000110;\
    conv2_weight_array[5][4][0][4] <= 18'b100000000010110100;\
    conv2_weight_array[5][4][1][0] <= 18'b100000000001011001;\
    conv2_weight_array[5][4][1][1] <= 18'b000000000010111100;\
    conv2_weight_array[5][4][1][2] <= 18'b000000000010000100;\
    conv2_weight_array[5][4][1][3] <= 18'b100000000011101011;\
    conv2_weight_array[5][4][1][4] <= 18'b100000000101010011;\
    conv2_weight_array[5][4][2][0] <= 18'b100000001001000011;\
    conv2_weight_array[5][4][2][1] <= 18'b100000000010000111;\
    conv2_weight_array[5][4][2][2] <= 18'b100000000000100101;\
    conv2_weight_array[5][4][2][3] <= 18'b000000000001010001;\
    conv2_weight_array[5][4][2][4] <= 18'b000000000000100110;\
    conv2_weight_array[5][4][3][0] <= 18'b000000000001011000;\
    conv2_weight_array[5][4][3][1] <= 18'b000000000010010011;\
    conv2_weight_array[5][4][3][2] <= 18'b000000000001101001;\
    conv2_weight_array[5][4][3][3] <= 18'b100000000011001100;\
    conv2_weight_array[5][4][3][4] <= 18'b100000000001111101;\
    conv2_weight_array[5][4][4][0] <= 18'b100000000000011110;\
    conv2_weight_array[5][4][4][1] <= 18'b100000000011011011;\
    conv2_weight_array[5][4][4][2] <= 18'b100000000010101001;\
    conv2_weight_array[5][4][4][3] <= 18'b100000000100010010;\
    conv2_weight_array[5][4][4][4] <= 18'b100000000010110011;\
    conv2_weight_array[5][5][0][0] <= 18'b100000000000100011;\
    conv2_weight_array[5][5][0][1] <= 18'b000000000000010011;\
    conv2_weight_array[5][5][0][2] <= 18'b000000000011101101;\
    conv2_weight_array[5][5][0][3] <= 18'b100000000100100011;\
    conv2_weight_array[5][5][0][4] <= 18'b100000000110001100;\
    conv2_weight_array[5][5][1][0] <= 18'b100000000000101011;\
    conv2_weight_array[5][5][1][1] <= 18'b100000000100001101;\
    conv2_weight_array[5][5][1][2] <= 18'b100000000000101111;\
    conv2_weight_array[5][5][1][3] <= 18'b000000000011001000;\
    conv2_weight_array[5][5][1][4] <= 18'b000000000110110010;\
    conv2_weight_array[5][5][2][0] <= 18'b100000000001011110;\
    conv2_weight_array[5][5][2][1] <= 18'b000000000001111110;\
    conv2_weight_array[5][5][2][2] <= 18'b000000000011100111;\
    conv2_weight_array[5][5][2][3] <= 18'b000000000101010111;\
    conv2_weight_array[5][5][2][4] <= 18'b000000000100101011;\
    conv2_weight_array[5][5][3][0] <= 18'b100000000100001110;\
    conv2_weight_array[5][5][3][1] <= 18'b100000000100000111;\
    conv2_weight_array[5][5][3][2] <= 18'b100000000101010110;\
    conv2_weight_array[5][5][3][3] <= 18'b000000000000000001;\
    conv2_weight_array[5][5][3][4] <= 18'b000000001000000101;\
    conv2_weight_array[5][5][4][0] <= 18'b100000000110100010;\
    conv2_weight_array[5][5][4][1] <= 18'b100000000001101000;\
    conv2_weight_array[5][5][4][2] <= 18'b100000000001110011;\
    conv2_weight_array[5][5][4][3] <= 18'b000000001100000100;\
    conv2_weight_array[5][5][4][4] <= 18'b000000001011100101;\
end