`define CACHE \
always@(posedge clk) begin\
    if((state>=CONV1_1_1)&(state<=CONV1_6_7)&(cnt2==8'd6))begin\
        cache[0] <= add_result[0];\
        cache[1] <= add_result[1];\
        cache[2] <= add_result[2];\
        cache[3] <= add_result[3];\
        cache[4] <= add_result[4];\
        cache[5] <= add_result[5];\
        cache[6] <= add_result[6];\
        cache[7] <= add_result[7];\
        cache[8] <= add_result[8];\
        cache[9] <= add_result[9];\
        cache[10] <= add_result[10];\
        cache[11] <= add_result[11];\
        cache[12] <= add_result[12];\
        cache[13] <= add_result[13];\
        cache[14] <= add_result[14];\
        cache[15] <= add_result[15];\
        cache[16] <= add_result[16];\
        cache[17] <= add_result[17];\
        cache[18] <= add_result[18];\
        cache[19] <= add_result[19];\
        cache[20] <= add_result[20];\
        cache[21] <= add_result[21];\
        cache[22] <= add_result[22];\
        cache[23] <= add_result[23];\
        cache[24] <= add_result[24];\
        cache[25] <= add_result[25];\
        cache[26] <= add_result[26];\
        cache[27] <= add_result[27];\
        cache[28] <= add_result[28];\
        cache[29] <= add_result[29];\
        cache[30] <= add_result[30];\
        cache[31] <= add_result[31];\
        cache[32] <= add_result[32];\
        cache[33] <= add_result[33];\
        cache[34] <= add_result[34];\
        cache[35] <= add_result[35];\
        cache[36] <= add_result[36];\
        cache[37] <= add_result[37];\
        cache[38] <= add_result[38];\
        cache[39] <= add_result[39];\
        cache[40] <= add_result[40];\
        cache[41] <= add_result[41];\
        cache[42] <= add_result[42];\
        cache[43] <= add_result[43];\
        cache[44] <= add_result[44];\
        cache[45] <= add_result[45];\
        cache[46] <= add_result[46];\
        cache[47] <= add_result[47];\
        cache[48] <= add_result[48];\
        cache[49] <= add_result[49];\
        cache[50] <= add_result[50];\
        cache[51] <= add_result[51];\
        cache[52] <= add_result[52];\
        cache[53] <= add_result[53];\
        cache[54] <= add_result[54];\
        cache[55] <= add_result[55];\
        cache[56] <= add_result[56];\
        cache[57] <= add_result[57];\
        cache[58] <= add_result[58];\
        cache[59] <= add_result[59];\
        cache[60] <= add_result[60];\
        cache[61] <= add_result[61];\
        cache[62] <= add_result[62];\
        cache[63] <= add_result[63];\
        cache[64] <= add_result[64];\
        cache[65] <= add_result[65];\
        cache[66] <= add_result[66];\
        cache[67] <= add_result[67];\
        cache[68] <= add_result[68];\
        cache[69] <= add_result[69];\
        cache[70] <= add_result[70];\
        cache[71] <= add_result[71];\
        cache[72] <= add_result[72];\
        cache[73] <= add_result[73];\
        cache[74] <= add_result[74];\
        cache[75] <= add_result[75];\
        cache[76] <= add_result[76];\
        cache[77] <= add_result[77];\
        cache[78] <= add_result[78];\
        cache[79] <= add_result[79];\
        cache[80] <= add_result[80];\
        cache[81] <= add_result[81];\
        cache[82] <= add_result[82];\
        cache[83] <= add_result[83];\
        cache[84] <= add_result[84];\
        cache[85] <= add_result[85];\
        cache[86] <= add_result[86];\
        cache[87] <= add_result[87];\
        cache[88] <= add_result[88];\
        cache[89] <= add_result[89];\
        cache[90] <= add_result[90];\
        cache[91] <= add_result[91];\
        cache[92] <= add_result[92];\
        cache[93] <= add_result[93];\
        cache[94] <= add_result[94];\
        cache[95] <= add_result[95];\
        cache[96] <= add_result[96];\
        cache[97] <= add_result[97];\
        cache[98] <= add_result[98];\
        cache[99] <= add_result[99];\
        cache[100] <= add_result[100];\
        cache[101] <= add_result[101];\
        cache[102] <= add_result[102];\
        cache[103] <= add_result[103];\
        cache[104] <= add_result[104];\
        cache[105] <= add_result[105];\
        cache[106] <= add_result[106];\
        cache[107] <= add_result[107];\
        cache[108] <= add_result[108];\
        cache[109] <= add_result[109];\
        cache[110] <= add_result[110];\
        cache[111] <= add_result[111];\
    end\
    else if((state==CONV2_1_6)|(state==CONV2_2_6)|(state==CONV2_3_6)|(state==CONV2_4_6)|(state==CONV2_5_6)|(state==CONV2_6_6))begin\
        cache[0] <= add_result[0];\
        cache[1] <= add_result[1];\
        cache[2] <= add_result[2];\
        cache[3] <= add_result[3];\
        cache[4] <= add_result[4];\
        cache[5] <= add_result[5];\
        cache[6] <= add_result[6];\
        cache[7] <= add_result[7];\
        cache[8] <= add_result[8];\
        cache[9] <= add_result[9];\
        cache[10] <= add_result[10];\
        cache[11] <= add_result[11];\
        cache[12] <= add_result[12];\
        cache[13] <= add_result[13];\
        cache[14] <= add_result[14];\
        cache[15] <= add_result[15];\
        cache[16] <= add_result[16];\
        cache[17] <= add_result[17];\
        cache[18] <= add_result[18];\
        cache[19] <= add_result[19];\
        cache[20] <= add_result[20];\
        cache[21] <= add_result[21];\
        cache[22] <= add_result[22];\
        cache[23] <= add_result[23];\
        cache[24] <= add_result[24];\
        cache[25] <= add_result[25];\
        cache[26] <= add_result[26];\
        cache[27] <= add_result[27];\
        cache[28] <= add_result[28];\
        cache[29] <= add_result[29];\
        cache[30] <= add_result[30];\
        cache[31] <= add_result[31];\
        cache[32] <= add_result[32];\
        cache[33] <= add_result[33];\
        cache[34] <= add_result[34];\
        cache[35] <= add_result[35];\
        cache[36] <= add_result[36];\
        cache[37] <= add_result[37];\
        cache[38] <= add_result[38];\
        cache[39] <= add_result[39];\
        cache[40] <= add_result[40];\
        cache[41] <= add_result[41];\
        cache[42] <= add_result[42];\
        cache[43] <= add_result[43];\
        cache[44] <= add_result[44];\
        cache[45] <= add_result[45];\
        cache[46] <= add_result[46];\
        cache[47] <= add_result[47];\
        cache[48] <= add_result[48];\
        cache[49] <= add_result[49];\
        cache[50] <= add_result[50];\
        cache[51] <= add_result[51];\
        cache[52] <= add_result[52];\
        cache[53] <= add_result[53];\
        cache[54] <= add_result[54];\
        cache[55] <= add_result[55];\
        cache[56] <= add_result[56];\
        cache[57] <= add_result[57];\
        cache[58] <= add_result[58];\
        cache[59] <= add_result[59];\
        cache[60] <= add_result[60];\
        cache[61] <= add_result[61];\
        cache[62] <= add_result[62];\
        cache[63] <= add_result[63];\
        cache[64] <= add_result[64];\
        cache[65] <= add_result[65];\
        cache[66] <= add_result[66];\
        cache[67] <= add_result[67];\
        cache[68] <= add_result[68];\
        cache[69] <= add_result[69];\
        cache[70] <= add_result[70];\
        cache[71] <= add_result[71];\
        cache[72] <= add_result[72];\
        cache[73] <= add_result[73];\
        cache[74] <= add_result[74];\
        cache[75] <= add_result[75];\
        cache[76] <= add_result[76];\
        cache[77] <= add_result[77];\
        cache[78] <= add_result[78];\
        cache[79] <= add_result[79];\
        cache[80] <= add_result[80];\
        cache[81] <= add_result[81];\
        cache[82] <= add_result[82];\
        cache[83] <= add_result[83];\
        cache[84] <= add_result[84];\
        cache[85] <= add_result[85];\
        cache[86] <= add_result[86];\
        cache[87] <= add_result[87];\
        cache[88] <= add_result[88];\
        cache[89] <= add_result[89];\
        cache[90] <= add_result[90];\
        cache[91] <= add_result[91];\
        cache[92] <= add_result[92];\
        cache[93] <= add_result[93];\
        cache[94] <= add_result[94];\
        cache[95] <= add_result[95];\
        cache[96] <= add_result[96];\
        cache[97] <= add_result[97];\
        cache[98] <= add_result[98];\
        cache[99] <= add_result[99];\
    end\
    else if(cnt1==8'd151) begin\
        cache[100] <= add_result[100][0] ? 18'd0 : add_result[100];\
        cache[101] <= add_result[101][0] ? 18'd0 : add_result[101];\
        cache[102] <= add_result[102][0] ? 18'd0 : add_result[102];\
        cache[103] <= add_result[103][0] ? 18'd0 : add_result[103];\
        cache[104] <= add_result[104][0] ? 18'd0 : add_result[104];\
        cache[105] <= add_result[105][0] ? 18'd0 : add_result[105];\
        cache[106] <= add_result[106][0] ? 18'd0 : add_result[106];\
        cache[107] <= add_result[107][0] ? 18'd0 : add_result[107];\
        cache[108] <= add_result[108][0] ? 18'd0 : add_result[108];\
        cache[109] <= add_result[109][0] ? 18'd0 : add_result[109];\
        cache[110] <= add_result[110][0] ? 18'd0 : add_result[110];\
        cache[111] <= add_result[111][0] ? 18'd0 : add_result[111];\
    end\
end