// `define CONV1_WEIGHT \
// reg [0:449] conv1_weight_array [0:5];\
// always@(posedge clk or negedge rst_n) begin\
//     conv1_weight_array[0] <= {25{18'h00400}};\
//     conv1_weight_array[1] <= {25{18'h00400}};\
//     conv1_weight_array[2] <= {25{18'h00400}};\
//     conv1_weight_array[3] <= {25{18'h00400}};\
//     conv1_weight_array[4] <= {25{18'h00400}};\
//     conv1_weight_array[5] <= {25{18'h00400}};\
// end

`define CONV1_WEIGHT \
reg [0:17] conv1_weight_array [0:5][0:4][0:4];\
always@(posedge clk) begin\
    conv1_weight_array[0][0][0] <= 18'b000000000101101100;\
    conv1_weight_array[0][0][1] <= 18'b100000000110011010;\
    conv1_weight_array[0][0][2] <= 18'b100000001101001011;\
    conv1_weight_array[0][0][3] <= 18'b100000000010100010;\
    conv1_weight_array[0][0][4] <= 18'b100000000000010001;\
    conv1_weight_array[0][1][0] <= 18'b000000001000000000;\
    conv1_weight_array[0][1][1] <= 18'b000000000000011010;\
    conv1_weight_array[0][1][2] <= 18'b100000001011111011;\
    conv1_weight_array[0][1][3] <= 18'b100000001010110100;\
    conv1_weight_array[0][1][4] <= 18'b100000001010101111;\
    conv1_weight_array[0][2][0] <= 18'b000000000101101101;\
    conv1_weight_array[0][2][1] <= 18'b000000000101101001;\
    conv1_weight_array[0][2][2] <= 18'b000000000000110111;\
    conv1_weight_array[0][2][3] <= 18'b000000000000000101;\
    conv1_weight_array[0][2][4] <= 18'b100000000011110001;\
    conv1_weight_array[0][3][0] <= 18'b000000000111100001;\
    conv1_weight_array[0][3][1] <= 18'b000000001010111001;\
    conv1_weight_array[0][3][2] <= 18'b000000000111111110;\
    conv1_weight_array[0][3][3] <= 18'b000000001000100111;\
    conv1_weight_array[0][3][4] <= 18'b000000000010001101;\
    conv1_weight_array[0][4][0] <= 18'b000000000010100001;\
    conv1_weight_array[0][4][1] <= 18'b000000000111000000;\
    conv1_weight_array[0][4][2] <= 18'b000000000111000001;\
    conv1_weight_array[0][4][3] <= 18'b000000000100011001;\
    conv1_weight_array[0][4][4] <= 18'b000000000110010000;\
    conv1_weight_array[1][0][0] <= 18'b000000000011110000;\
    conv1_weight_array[1][0][1] <= 18'b100000000101001010;\
    conv1_weight_array[1][0][2] <= 18'b100000000101101110;\
    conv1_weight_array[1][0][3] <= 18'b000000000000100111;\
    conv1_weight_array[1][0][4] <= 18'b000000000111010000;\
    conv1_weight_array[1][1][0] <= 18'b100000000110101001;\
    conv1_weight_array[1][1][1] <= 18'b100000000011111100;\
    conv1_weight_array[1][1][2] <= 18'b000000000110001000;\
    conv1_weight_array[1][1][3] <= 18'b000000001000001001;\
    conv1_weight_array[1][1][4] <= 18'b000000000101000111;\
    conv1_weight_array[1][2][0] <= 18'b100000000001100111;\
    conv1_weight_array[1][2][1] <= 18'b000000000110100001;\
    conv1_weight_array[1][2][2] <= 18'b000000001110011011;\
    conv1_weight_array[1][2][3] <= 18'b000000001101000110;\
    conv1_weight_array[1][2][4] <= 18'b100000000000100110;\
    conv1_weight_array[1][3][0] <= 18'b100000000011000111;\
    conv1_weight_array[1][3][1] <= 18'b000000000011010110;\
    conv1_weight_array[1][3][2] <= 18'b000000000100101110;\
    conv1_weight_array[1][3][3] <= 18'b100000000101010001;\
    conv1_weight_array[1][3][4] <= 18'b100000001111011001;\
    conv1_weight_array[1][4][0] <= 18'b000000000010011100;\
    conv1_weight_array[1][4][1] <= 18'b000000000011100001;\
    conv1_weight_array[1][4][2] <= 18'b100000000110100101;\
    conv1_weight_array[1][4][3] <= 18'b100000001101111110;\
    conv1_weight_array[1][4][4] <= 18'b100000001001100110;\
    conv1_weight_array[2][0][0] <= 18'b100000000001001110;\
    conv1_weight_array[2][0][1] <= 18'b000000000101010010;\
    conv1_weight_array[2][0][2] <= 18'b000000000011111000;\
    conv1_weight_array[2][0][3] <= 18'b100000000101011000;\
    conv1_weight_array[2][0][4] <= 18'b100000000000010001;\
    conv1_weight_array[2][1][0] <= 18'b100000000001100100;\
    conv1_weight_array[2][1][1] <= 18'b000000000111101011;\
    conv1_weight_array[2][1][2] <= 18'b000000000000011111;\
    conv1_weight_array[2][1][3] <= 18'b100000001001011000;\
    conv1_weight_array[2][1][4] <= 18'b000000000010101100;\
    conv1_weight_array[2][2][0] <= 18'b000000000011101011;\
    conv1_weight_array[2][2][1] <= 18'b000000001011000110;\
    conv1_weight_array[2][2][2] <= 18'b100000000100010101;\
    conv1_weight_array[2][2][3] <= 18'b000000000001100101;\
    conv1_weight_array[2][2][4] <= 18'b000000001000101111;\
    conv1_weight_array[2][3][0] <= 18'b100000000000100111;\
    conv1_weight_array[2][3][1] <= 18'b000000001001001000;\
    conv1_weight_array[2][3][2] <= 18'b000000000010001011;\
    conv1_weight_array[2][3][3] <= 18'b000000000001011101;\
    conv1_weight_array[2][3][4] <= 18'b000000001001000011;\
    conv1_weight_array[2][4][0] <= 18'b100000000010101001;\
    conv1_weight_array[2][4][1] <= 18'b000000000100111011;\
    conv1_weight_array[2][4][2] <= 18'b100000000000001011;\
    conv1_weight_array[2][4][3] <= 18'b100000000101011111;\
    conv1_weight_array[2][4][4] <= 18'b100000000000001010;\
    conv1_weight_array[3][0][0] <= 18'b100000000011011010;\
    conv1_weight_array[3][0][1] <= 18'b000000000001101011;\
    conv1_weight_array[3][0][2] <= 18'b000000000110001111;\
    conv1_weight_array[3][0][3] <= 18'b000000000011100001;\
    conv1_weight_array[3][0][4] <= 18'b000000000010100000;\
    conv1_weight_array[3][1][0] <= 18'b100000000000010000;\
    conv1_weight_array[3][1][1] <= 18'b000000000100100111;\
    conv1_weight_array[3][1][2] <= 18'b000000000111111110;\
    conv1_weight_array[3][1][3] <= 18'b000000000000000010;\
    conv1_weight_array[3][1][4] <= 18'b100000000000010101;\
    conv1_weight_array[3][2][0] <= 18'b100000000000011100;\
    conv1_weight_array[3][2][1] <= 18'b000000000101111011;\
    conv1_weight_array[3][2][2] <= 18'b000000000111110011;\
    conv1_weight_array[3][2][3] <= 18'b000000000001011011;\
    conv1_weight_array[3][2][4] <= 18'b000000000001100101;\
    conv1_weight_array[3][3][0] <= 18'b000000000011010100;\
    conv1_weight_array[3][3][1] <= 18'b000000000110101101;\
    conv1_weight_array[3][3][2] <= 18'b000000000111010010;\
    conv1_weight_array[3][3][3] <= 18'b100000000000011011;\
    conv1_weight_array[3][3][4] <= 18'b000000000001001101;\
    conv1_weight_array[3][4][0] <= 18'b000000000010000011;\
    conv1_weight_array[3][4][1] <= 18'b000000000011101000;\
    conv1_weight_array[3][4][2] <= 18'b000000001000110100;\
    conv1_weight_array[3][4][3] <= 18'b000000000100101011;\
    conv1_weight_array[3][4][4] <= 18'b000000000011000101;\
    conv1_weight_array[4][0][0] <= 18'b000000000100001110;\
    conv1_weight_array[4][0][1] <= 18'b000000000110100101;\
    conv1_weight_array[4][0][2] <= 18'b000000000111000010;\
    conv1_weight_array[4][0][3] <= 18'b100000000011100000;\
    conv1_weight_array[4][0][4] <= 18'b100000010000111000;\
    conv1_weight_array[4][1][0] <= 18'b000000000011001110;\
    conv1_weight_array[4][1][1] <= 18'b000000000101011011;\
    conv1_weight_array[4][1][2] <= 18'b000000000001100000;\
    conv1_weight_array[4][1][3] <= 18'b100000000101100111;\
    conv1_weight_array[4][1][4] <= 18'b100000010101011110;\
    conv1_weight_array[4][2][0] <= 18'b000000001000111111;\
    conv1_weight_array[4][2][1] <= 18'b000000000100100100;\
    conv1_weight_array[4][2][2] <= 18'b100000000000100101;\
    conv1_weight_array[4][2][3] <= 18'b100000001011110101;\
    conv1_weight_array[4][2][4] <= 18'b100000010100010000;\
    conv1_weight_array[4][3][0] <= 18'b000000000111010101;\
    conv1_weight_array[4][3][1] <= 18'b000000000010111011;\
    conv1_weight_array[4][3][2] <= 18'b100000000010100001;\
    conv1_weight_array[4][3][3] <= 18'b100000001111101101;\
    conv1_weight_array[4][3][4] <= 18'b100000001001001010;\
    conv1_weight_array[4][4][0] <= 18'b000000001000100111;\
    conv1_weight_array[4][4][1] <= 18'b000000000011011001;\
    conv1_weight_array[4][4][2] <= 18'b100000001010000011;\
    conv1_weight_array[4][4][3] <= 18'b100000001111001000;\
    conv1_weight_array[4][4][4] <= 18'b000000000000111010;\
    conv1_weight_array[5][0][0] <= 18'b000000000001101100;\
    conv1_weight_array[5][0][1] <= 18'b000000000001101111;\
    conv1_weight_array[5][0][2] <= 18'b000000000011111100;\
    conv1_weight_array[5][0][3] <= 18'b100000000000110010;\
    conv1_weight_array[5][0][4] <= 18'b100000000100000110;\
    conv1_weight_array[5][1][0] <= 18'b000000001010001010;\
    conv1_weight_array[5][1][1] <= 18'b000000000101111110;\
    conv1_weight_array[5][1][2] <= 18'b000000000100100001;\
    conv1_weight_array[5][1][3] <= 18'b100000000111000010;\
    conv1_weight_array[5][1][4] <= 18'b100000000101010011;\
    conv1_weight_array[5][2][0] <= 18'b000000000010100000;\
    conv1_weight_array[5][2][1] <= 18'b100000001000101111;\
    conv1_weight_array[5][2][2] <= 18'b100000001011011110;\
    conv1_weight_array[5][2][3] <= 18'b100000001100000010;\
    conv1_weight_array[5][2][4] <= 18'b000000000011010110;\
    conv1_weight_array[5][3][0] <= 18'b100000000011010001;\
    conv1_weight_array[5][3][1] <= 18'b100000001100000011;\
    conv1_weight_array[5][3][2] <= 18'b100000000110110011;\
    conv1_weight_array[5][3][3] <= 18'b000000001000011101;\
    conv1_weight_array[5][3][4] <= 18'b000000001011111110;\
    conv1_weight_array[5][4][0] <= 18'b100000000000011010;\
    conv1_weight_array[5][4][1] <= 18'b000000000011100010;\
    conv1_weight_array[5][4][2] <= 18'b000000000101110101;\
    conv1_weight_array[5][4][3] <= 18'b000000000110011000;\
    conv1_weight_array[5][4][4] <= 18'b100000000001010011;\
end