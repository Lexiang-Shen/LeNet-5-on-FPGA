`define IN_IMG_ARRAY \
always@(posedge clk or negedge rst_n) begin\
    if(!rst_n) begin\
        in_img_array[0][0] <= 18'd0;\
        in_img_array[0][1] <= 18'd0;\
        in_img_array[0][2] <= 18'd0;\
        in_img_array[0][3] <= 18'd0;\
        in_img_array[0][4] <= 18'd0;\
        in_img_array[0][5] <= 18'd0;\
        in_img_array[0][6] <= 18'd0;\
        in_img_array[0][7] <= 18'd0;\
        in_img_array[0][8] <= 18'd0;\
        in_img_array[0][9] <= 18'd0;\
        in_img_array[0][10] <= 18'd0;\
        in_img_array[0][11] <= 18'd0;\
        in_img_array[0][12] <= 18'd0;\
        in_img_array[0][13] <= 18'd0;\
        in_img_array[0][14] <= 18'd0;\
        in_img_array[0][15] <= 18'd0;\
        in_img_array[0][16] <= 18'd0;\
        in_img_array[0][17] <= 18'd0;\
        in_img_array[0][18] <= 18'd0;\
        in_img_array[0][19] <= 18'd0;\
        in_img_array[0][20] <= 18'd0;\
        in_img_array[0][21] <= 18'd0;\
        in_img_array[0][22] <= 18'd0;\
        in_img_array[0][23] <= 18'd0;\
        in_img_array[0][24] <= 18'd0;\
        in_img_array[0][25] <= 18'd0;\
        in_img_array[0][26] <= 18'd0;\
        in_img_array[0][27] <= 18'd0;\
        in_img_array[0][28] <= 18'd0;\
        in_img_array[0][29] <= 18'd0;\
        in_img_array[0][30] <= 18'd0;\
        in_img_array[0][31] <= 18'd0;\
        in_img_array[1][0] <= 18'd0;\
        in_img_array[1][1] <= 18'd0;\
        in_img_array[1][2] <= 18'd0;\
        in_img_array[1][3] <= 18'd0;\
        in_img_array[1][4] <= 18'd0;\
        in_img_array[1][5] <= 18'd0;\
        in_img_array[1][6] <= 18'd0;\
        in_img_array[1][7] <= 18'd0;\
        in_img_array[1][8] <= 18'd0;\
        in_img_array[1][9] <= 18'd0;\
        in_img_array[1][10] <= 18'd0;\
        in_img_array[1][11] <= 18'd0;\
        in_img_array[1][12] <= 18'd0;\
        in_img_array[1][13] <= 18'd0;\
        in_img_array[1][14] <= 18'd0;\
        in_img_array[1][15] <= 18'd0;\
        in_img_array[1][16] <= 18'd0;\
        in_img_array[1][17] <= 18'd0;\
        in_img_array[1][18] <= 18'd0;\
        in_img_array[1][19] <= 18'd0;\
        in_img_array[1][20] <= 18'd0;\
        in_img_array[1][21] <= 18'd0;\
        in_img_array[1][22] <= 18'd0;\
        in_img_array[1][23] <= 18'd0;\
        in_img_array[1][24] <= 18'd0;\
        in_img_array[1][25] <= 18'd0;\
        in_img_array[1][26] <= 18'd0;\
        in_img_array[1][27] <= 18'd0;\
        in_img_array[1][28] <= 18'd0;\
        in_img_array[1][29] <= 18'd0;\
        in_img_array[1][30] <= 18'd0;\
        in_img_array[1][31] <= 18'd0;\
        in_img_array[2][0] <= 18'd0;\
        in_img_array[2][1] <= 18'd0;\
        in_img_array[2][2] <= 18'd0;\
        in_img_array[2][3] <= 18'd0;\
        in_img_array[2][4] <= 18'd0;\
        in_img_array[2][5] <= 18'd0;\
        in_img_array[2][6] <= 18'd0;\
        in_img_array[2][7] <= 18'd0;\
        in_img_array[2][8] <= 18'd0;\
        in_img_array[2][9] <= 18'd0;\
        in_img_array[2][10] <= 18'd0;\
        in_img_array[2][11] <= 18'd0;\
        in_img_array[2][12] <= 18'd0;\
        in_img_array[2][13] <= 18'd0;\
        in_img_array[2][14] <= 18'd0;\
        in_img_array[2][15] <= 18'd0;\
        in_img_array[2][16] <= 18'd0;\
        in_img_array[2][17] <= 18'd0;\
        in_img_array[2][18] <= 18'd0;\
        in_img_array[2][19] <= 18'd0;\
        in_img_array[2][20] <= 18'd0;\
        in_img_array[2][21] <= 18'd0;\
        in_img_array[2][22] <= 18'd0;\
        in_img_array[2][23] <= 18'd0;\
        in_img_array[2][24] <= 18'd0;\
        in_img_array[2][25] <= 18'd0;\
        in_img_array[2][26] <= 18'd0;\
        in_img_array[2][27] <= 18'd0;\
        in_img_array[2][28] <= 18'd0;\
        in_img_array[2][29] <= 18'd0;\
        in_img_array[2][30] <= 18'd0;\
        in_img_array[2][31] <= 18'd0;\
        in_img_array[3][0] <= 18'd0;\
        in_img_array[3][1] <= 18'd0;\
        in_img_array[3][2] <= 18'd0;\
        in_img_array[3][3] <= 18'd0;\
        in_img_array[3][4] <= 18'd0;\
        in_img_array[3][5] <= 18'd0;\
        in_img_array[3][6] <= 18'd0;\
        in_img_array[3][7] <= 18'd0;\
        in_img_array[3][8] <= 18'd0;\
        in_img_array[3][9] <= 18'd0;\
        in_img_array[3][10] <= 18'd0;\
        in_img_array[3][11] <= 18'd0;\
        in_img_array[3][12] <= 18'd0;\
        in_img_array[3][13] <= 18'd0;\
        in_img_array[3][14] <= 18'd0;\
        in_img_array[3][15] <= 18'd0;\
        in_img_array[3][16] <= 18'd0;\
        in_img_array[3][17] <= 18'd0;\
        in_img_array[3][18] <= 18'd0;\
        in_img_array[3][19] <= 18'd0;\
        in_img_array[3][20] <= 18'd0;\
        in_img_array[3][21] <= 18'd0;\
        in_img_array[3][22] <= 18'd0;\
        in_img_array[3][23] <= 18'd0;\
        in_img_array[3][24] <= 18'd0;\
        in_img_array[3][25] <= 18'd0;\
        in_img_array[3][26] <= 18'd0;\
        in_img_array[3][27] <= 18'd0;\
        in_img_array[3][28] <= 18'd0;\
        in_img_array[3][29] <= 18'd0;\
        in_img_array[3][30] <= 18'd0;\
        in_img_array[3][31] <= 18'd0;\
        in_img_array[4][0] <= 18'd0;\
        in_img_array[4][1] <= 18'd0;\
        in_img_array[4][2] <= 18'd0;\
        in_img_array[4][3] <= 18'd0;\
        in_img_array[4][4] <= 18'd0;\
        in_img_array[4][5] <= 18'd0;\
        in_img_array[4][6] <= 18'd0;\
        in_img_array[4][7] <= 18'd0;\
        in_img_array[4][8] <= 18'd0;\
        in_img_array[4][9] <= 18'd0;\
        in_img_array[4][10] <= 18'd0;\
        in_img_array[4][11] <= 18'd0;\
        in_img_array[4][12] <= 18'd0;\
        in_img_array[4][13] <= 18'd0;\
        in_img_array[4][14] <= 18'd0;\
        in_img_array[4][15] <= 18'd0;\
        in_img_array[4][16] <= 18'd0;\
        in_img_array[4][17] <= 18'd0;\
        in_img_array[4][18] <= 18'd0;\
        in_img_array[4][19] <= 18'd0;\
        in_img_array[4][20] <= 18'd0;\
        in_img_array[4][21] <= 18'd0;\
        in_img_array[4][22] <= 18'd0;\
        in_img_array[4][23] <= 18'd0;\
        in_img_array[4][24] <= 18'd0;\
        in_img_array[4][25] <= 18'd0;\
        in_img_array[4][26] <= 18'd0;\
        in_img_array[4][27] <= 18'd0;\
        in_img_array[4][28] <= 18'd0;\
        in_img_array[4][29] <= 18'd0;\
        in_img_array[4][30] <= 18'd0;\
        in_img_array[4][31] <= 18'd0;\
        in_img_array[5][0] <= 18'd0;\
        in_img_array[5][1] <= 18'd0;\
        in_img_array[5][2] <= 18'd0;\
        in_img_array[5][3] <= 18'd0;\
        in_img_array[5][4] <= 18'd0;\
        in_img_array[5][5] <= 18'd0;\
        in_img_array[5][6] <= 18'd0;\
        in_img_array[5][7] <= 18'd0;\
        in_img_array[5][8] <= 18'd0;\
        in_img_array[5][9] <= 18'd0;\
        in_img_array[5][10] <= 18'd0;\
        in_img_array[5][11] <= 18'd0;\
        in_img_array[5][12] <= 18'd0;\
        in_img_array[5][13] <= 18'd0;\
        in_img_array[5][14] <= 18'd0;\
        in_img_array[5][15] <= 18'd0;\
        in_img_array[5][16] <= 18'd0;\
        in_img_array[5][17] <= 18'd0;\
        in_img_array[5][18] <= 18'd0;\
        in_img_array[5][19] <= 18'd0;\
        in_img_array[5][20] <= 18'd0;\
        in_img_array[5][21] <= 18'd0;\
        in_img_array[5][22] <= 18'd0;\
        in_img_array[5][23] <= 18'd0;\
        in_img_array[5][24] <= 18'd0;\
        in_img_array[5][25] <= 18'd0;\
        in_img_array[5][26] <= 18'd0;\
        in_img_array[5][27] <= 18'd0;\
        in_img_array[5][28] <= 18'd0;\
        in_img_array[5][29] <= 18'd0;\
        in_img_array[5][30] <= 18'd0;\
        in_img_array[5][31] <= 18'd0;\
        in_img_array[6][0] <= 18'd0;\
        in_img_array[6][1] <= 18'd0;\
        in_img_array[6][2] <= 18'd0;\
        in_img_array[6][3] <= 18'd0;\
        in_img_array[6][4] <= 18'd0;\
        in_img_array[6][5] <= 18'd0;\
        in_img_array[6][6] <= 18'd0;\
        in_img_array[6][7] <= 18'd0;\
        in_img_array[6][8] <= 18'd0;\
        in_img_array[6][9] <= 18'd0;\
        in_img_array[6][10] <= 18'd0;\
        in_img_array[6][11] <= 18'd0;\
        in_img_array[6][12] <= 18'd0;\
        in_img_array[6][13] <= 18'd0;\
        in_img_array[6][14] <= 18'd0;\
        in_img_array[6][15] <= 18'd0;\
        in_img_array[6][16] <= 18'd0;\
        in_img_array[6][17] <= 18'd0;\
        in_img_array[6][18] <= 18'd0;\
        in_img_array[6][19] <= 18'd0;\
        in_img_array[6][20] <= 18'd0;\
        in_img_array[6][21] <= 18'd0;\
        in_img_array[6][22] <= 18'd0;\
        in_img_array[6][23] <= 18'd0;\
        in_img_array[6][24] <= 18'd0;\
        in_img_array[6][25] <= 18'd0;\
        in_img_array[6][26] <= 18'd0;\
        in_img_array[6][27] <= 18'd0;\
        in_img_array[6][28] <= 18'd0;\
        in_img_array[6][29] <= 18'd0;\
        in_img_array[6][30] <= 18'd0;\
        in_img_array[6][31] <= 18'd0;\
        in_img_array[7][0] <= 18'd0;\
        in_img_array[7][1] <= 18'd0;\
        in_img_array[7][2] <= 18'd0;\
        in_img_array[7][3] <= 18'd0;\
        in_img_array[7][4] <= 18'd0;\
        in_img_array[7][5] <= 18'd0;\
        in_img_array[7][6] <= 18'd0;\
        in_img_array[7][7] <= 18'd0;\
        in_img_array[7][8] <= 18'd0;\
        in_img_array[7][9] <= 18'd0;\
        in_img_array[7][10] <= 18'd0;\
        in_img_array[7][11] <= 18'd0;\
        in_img_array[7][12] <= 18'd0;\
        in_img_array[7][13] <= 18'd0;\
        in_img_array[7][14] <= 18'd0;\
        in_img_array[7][15] <= 18'd0;\
        in_img_array[7][16] <= 18'd0;\
        in_img_array[7][17] <= 18'd0;\
        in_img_array[7][18] <= 18'd0;\
        in_img_array[7][19] <= 18'd0;\
        in_img_array[7][20] <= 18'd0;\
        in_img_array[7][21] <= 18'd0;\
        in_img_array[7][22] <= 18'd0;\
        in_img_array[7][23] <= 18'd0;\
        in_img_array[7][24] <= 18'd0;\
        in_img_array[7][25] <= 18'd0;\
        in_img_array[7][26] <= 18'd0;\
        in_img_array[7][27] <= 18'd0;\
        in_img_array[7][28] <= 18'd0;\
        in_img_array[7][29] <= 18'd0;\
        in_img_array[7][30] <= 18'd0;\
        in_img_array[7][31] <= 18'd0;\
        in_img_array[8][0] <= 18'd0;\
        in_img_array[8][1] <= 18'd0;\
        in_img_array[8][2] <= 18'd0;\
        in_img_array[8][3] <= 18'd0;\
        in_img_array[8][4] <= 18'd0;\
        in_img_array[8][5] <= 18'd0;\
        in_img_array[8][6] <= 18'd0;\
        in_img_array[8][7] <= 18'd0;\
        in_img_array[8][8] <= 18'd0;\
        in_img_array[8][9] <= 18'd0;\
        in_img_array[8][10] <= 18'd0;\
        in_img_array[8][11] <= 18'd0;\
        in_img_array[8][12] <= 18'd0;\
        in_img_array[8][13] <= 18'd0;\
        in_img_array[8][14] <= 18'd0;\
        in_img_array[8][15] <= 18'd0;\
        in_img_array[8][16] <= 18'd0;\
        in_img_array[8][17] <= 18'd0;\
        in_img_array[8][18] <= 18'd0;\
        in_img_array[8][19] <= 18'd0;\
        in_img_array[8][20] <= 18'd0;\
        in_img_array[8][21] <= 18'd0;\
        in_img_array[8][22] <= 18'd0;\
        in_img_array[8][23] <= 18'd0;\
        in_img_array[8][24] <= 18'd0;\
        in_img_array[8][25] <= 18'd0;\
        in_img_array[8][26] <= 18'd0;\
        in_img_array[8][27] <= 18'd0;\
        in_img_array[8][28] <= 18'd0;\
        in_img_array[8][29] <= 18'd0;\
        in_img_array[8][30] <= 18'd0;\
        in_img_array[8][31] <= 18'd0;\
        in_img_array[9][0] <= 18'd0;\
        in_img_array[9][1] <= 18'd0;\
        in_img_array[9][2] <= 18'd0;\
        in_img_array[9][3] <= 18'd0;\
        in_img_array[9][4] <= 18'd0;\
        in_img_array[9][5] <= 18'd0;\
        in_img_array[9][6] <= 18'd0;\
        in_img_array[9][7] <= 18'd0;\
        in_img_array[9][8] <= 18'd0;\
        in_img_array[9][9] <= 18'd0;\
        in_img_array[9][10] <= 18'd0;\
        in_img_array[9][11] <= 18'd0;\
        in_img_array[9][12] <= 18'd0;\
        in_img_array[9][13] <= 18'd0;\
        in_img_array[9][14] <= 18'd0;\
        in_img_array[9][15] <= 18'd0;\
        in_img_array[9][16] <= 18'd0;\
        in_img_array[9][17] <= 18'd0;\
        in_img_array[9][18] <= 18'd0;\
        in_img_array[9][19] <= 18'd0;\
        in_img_array[9][20] <= 18'd0;\
        in_img_array[9][21] <= 18'd0;\
        in_img_array[9][22] <= 18'd0;\
        in_img_array[9][23] <= 18'd0;\
        in_img_array[9][24] <= 18'd0;\
        in_img_array[9][25] <= 18'd0;\
        in_img_array[9][26] <= 18'd0;\
        in_img_array[9][27] <= 18'd0;\
        in_img_array[9][28] <= 18'd0;\
        in_img_array[9][29] <= 18'd0;\
        in_img_array[9][30] <= 18'd0;\
        in_img_array[9][31] <= 18'd0;\
        in_img_array[10][0] <= 18'd0;\
        in_img_array[10][1] <= 18'd0;\
        in_img_array[10][2] <= 18'd0;\
        in_img_array[10][3] <= 18'd0;\
        in_img_array[10][4] <= 18'd0;\
        in_img_array[10][5] <= 18'd0;\
        in_img_array[10][6] <= 18'd0;\
        in_img_array[10][7] <= 18'd0;\
        in_img_array[10][8] <= 18'd0;\
        in_img_array[10][9] <= 18'd0;\
        in_img_array[10][10] <= 18'd0;\
        in_img_array[10][11] <= 18'd0;\
        in_img_array[10][12] <= 18'd0;\
        in_img_array[10][13] <= 18'd0;\
        in_img_array[10][14] <= 18'd0;\
        in_img_array[10][15] <= 18'd0;\
        in_img_array[10][16] <= 18'd0;\
        in_img_array[10][17] <= 18'd0;\
        in_img_array[10][18] <= 18'd0;\
        in_img_array[10][19] <= 18'd0;\
        in_img_array[10][20] <= 18'd0;\
        in_img_array[10][21] <= 18'd0;\
        in_img_array[10][22] <= 18'd0;\
        in_img_array[10][23] <= 18'd0;\
        in_img_array[10][24] <= 18'd0;\
        in_img_array[10][25] <= 18'd0;\
        in_img_array[10][26] <= 18'd0;\
        in_img_array[10][27] <= 18'd0;\
        in_img_array[10][28] <= 18'd0;\
        in_img_array[10][29] <= 18'd0;\
        in_img_array[10][30] <= 18'd0;\
        in_img_array[10][31] <= 18'd0;\
        in_img_array[11][0] <= 18'd0;\
        in_img_array[11][1] <= 18'd0;\
        in_img_array[11][2] <= 18'd0;\
        in_img_array[11][3] <= 18'd0;\
        in_img_array[11][4] <= 18'd0;\
        in_img_array[11][5] <= 18'd0;\
        in_img_array[11][6] <= 18'd0;\
        in_img_array[11][7] <= 18'd0;\
        in_img_array[11][8] <= 18'd0;\
        in_img_array[11][9] <= 18'd0;\
        in_img_array[11][10] <= 18'd0;\
        in_img_array[11][11] <= 18'd0;\
        in_img_array[11][12] <= 18'd0;\
        in_img_array[11][13] <= 18'd0;\
        in_img_array[11][14] <= 18'd0;\
        in_img_array[11][15] <= 18'd0;\
        in_img_array[11][16] <= 18'd0;\
        in_img_array[11][17] <= 18'd0;\
        in_img_array[11][18] <= 18'd0;\
        in_img_array[11][19] <= 18'd0;\
        in_img_array[11][20] <= 18'd0;\
        in_img_array[11][21] <= 18'd0;\
        in_img_array[11][22] <= 18'd0;\
        in_img_array[11][23] <= 18'd0;\
        in_img_array[11][24] <= 18'd0;\
        in_img_array[11][25] <= 18'd0;\
        in_img_array[11][26] <= 18'd0;\
        in_img_array[11][27] <= 18'd0;\
        in_img_array[11][28] <= 18'd0;\
        in_img_array[11][29] <= 18'd0;\
        in_img_array[11][30] <= 18'd0;\
        in_img_array[11][31] <= 18'd0;\
        in_img_array[12][0] <= 18'd0;\
        in_img_array[12][1] <= 18'd0;\
        in_img_array[12][2] <= 18'd0;\
        in_img_array[12][3] <= 18'd0;\
        in_img_array[12][4] <= 18'd0;\
        in_img_array[12][5] <= 18'd0;\
        in_img_array[12][6] <= 18'd0;\
        in_img_array[12][7] <= 18'd0;\
        in_img_array[12][8] <= 18'd0;\
        in_img_array[12][9] <= 18'd0;\
        in_img_array[12][10] <= 18'd0;\
        in_img_array[12][11] <= 18'd0;\
        in_img_array[12][12] <= 18'd0;\
        in_img_array[12][13] <= 18'd0;\
        in_img_array[12][14] <= 18'd0;\
        in_img_array[12][15] <= 18'd0;\
        in_img_array[12][16] <= 18'd0;\
        in_img_array[12][17] <= 18'd0;\
        in_img_array[12][18] <= 18'd0;\
        in_img_array[12][19] <= 18'd0;\
        in_img_array[12][20] <= 18'd0;\
        in_img_array[12][21] <= 18'd0;\
        in_img_array[12][22] <= 18'd0;\
        in_img_array[12][23] <= 18'd0;\
        in_img_array[12][24] <= 18'd0;\
        in_img_array[12][25] <= 18'd0;\
        in_img_array[12][26] <= 18'd0;\
        in_img_array[12][27] <= 18'd0;\
        in_img_array[12][28] <= 18'd0;\
        in_img_array[12][29] <= 18'd0;\
        in_img_array[12][30] <= 18'd0;\
        in_img_array[12][31] <= 18'd0;\
        in_img_array[13][0] <= 18'd0;\
        in_img_array[13][1] <= 18'd0;\
        in_img_array[13][2] <= 18'd0;\
        in_img_array[13][3] <= 18'd0;\
        in_img_array[13][4] <= 18'd0;\
        in_img_array[13][5] <= 18'd0;\
        in_img_array[13][6] <= 18'd0;\
        in_img_array[13][7] <= 18'd0;\
        in_img_array[13][8] <= 18'd0;\
        in_img_array[13][9] <= 18'd0;\
        in_img_array[13][10] <= 18'd0;\
        in_img_array[13][11] <= 18'd0;\
        in_img_array[13][12] <= 18'd0;\
        in_img_array[13][13] <= 18'd0;\
        in_img_array[13][14] <= 18'd0;\
        in_img_array[13][15] <= 18'd0;\
        in_img_array[13][16] <= 18'd0;\
        in_img_array[13][17] <= 18'd0;\
        in_img_array[13][18] <= 18'd0;\
        in_img_array[13][19] <= 18'd0;\
        in_img_array[13][20] <= 18'd0;\
        in_img_array[13][21] <= 18'd0;\
        in_img_array[13][22] <= 18'd0;\
        in_img_array[13][23] <= 18'd0;\
        in_img_array[13][24] <= 18'd0;\
        in_img_array[13][25] <= 18'd0;\
        in_img_array[13][26] <= 18'd0;\
        in_img_array[13][27] <= 18'd0;\
        in_img_array[13][28] <= 18'd0;\
        in_img_array[13][29] <= 18'd0;\
        in_img_array[13][30] <= 18'd0;\
        in_img_array[13][31] <= 18'd0;\
        in_img_array[14][0] <= 18'd0;\
        in_img_array[14][1] <= 18'd0;\
        in_img_array[14][2] <= 18'd0;\
        in_img_array[14][3] <= 18'd0;\
        in_img_array[14][4] <= 18'd0;\
        in_img_array[14][5] <= 18'd0;\
        in_img_array[14][6] <= 18'd0;\
        in_img_array[14][7] <= 18'd0;\
        in_img_array[14][8] <= 18'd0;\
        in_img_array[14][9] <= 18'd0;\
        in_img_array[14][10] <= 18'd0;\
        in_img_array[14][11] <= 18'd0;\
        in_img_array[14][12] <= 18'd0;\
        in_img_array[14][13] <= 18'd0;\
        in_img_array[14][14] <= 18'd0;\
        in_img_array[14][15] <= 18'd0;\
        in_img_array[14][16] <= 18'd0;\
        in_img_array[14][17] <= 18'd0;\
        in_img_array[14][18] <= 18'd0;\
        in_img_array[14][19] <= 18'd0;\
        in_img_array[14][20] <= 18'd0;\
        in_img_array[14][21] <= 18'd0;\
        in_img_array[14][22] <= 18'd0;\
        in_img_array[14][23] <= 18'd0;\
        in_img_array[14][24] <= 18'd0;\
        in_img_array[14][25] <= 18'd0;\
        in_img_array[14][26] <= 18'd0;\
        in_img_array[14][27] <= 18'd0;\
        in_img_array[14][28] <= 18'd0;\
        in_img_array[14][29] <= 18'd0;\
        in_img_array[14][30] <= 18'd0;\
        in_img_array[14][31] <= 18'd0;\
        in_img_array[15][0] <= 18'd0;\
        in_img_array[15][1] <= 18'd0;\
        in_img_array[15][2] <= 18'd0;\
        in_img_array[15][3] <= 18'd0;\
        in_img_array[15][4] <= 18'd0;\
        in_img_array[15][5] <= 18'd0;\
        in_img_array[15][6] <= 18'd0;\
        in_img_array[15][7] <= 18'd0;\
        in_img_array[15][8] <= 18'd0;\
        in_img_array[15][9] <= 18'd0;\
        in_img_array[15][10] <= 18'd0;\
        in_img_array[15][11] <= 18'd0;\
        in_img_array[15][12] <= 18'd0;\
        in_img_array[15][13] <= 18'd0;\
        in_img_array[15][14] <= 18'd0;\
        in_img_array[15][15] <= 18'd0;\
        in_img_array[15][16] <= 18'd0;\
        in_img_array[15][17] <= 18'd0;\
        in_img_array[15][18] <= 18'd0;\
        in_img_array[15][19] <= 18'd0;\
        in_img_array[15][20] <= 18'd0;\
        in_img_array[15][21] <= 18'd0;\
        in_img_array[15][22] <= 18'd0;\
        in_img_array[15][23] <= 18'd0;\
        in_img_array[15][24] <= 18'd0;\
        in_img_array[15][25] <= 18'd0;\
        in_img_array[15][26] <= 18'd0;\
        in_img_array[15][27] <= 18'd0;\
        in_img_array[15][28] <= 18'd0;\
        in_img_array[15][29] <= 18'd0;\
        in_img_array[15][30] <= 18'd0;\
        in_img_array[15][31] <= 18'd0;\
        in_img_array[16][0] <= 18'd0;\
        in_img_array[16][1] <= 18'd0;\
        in_img_array[16][2] <= 18'd0;\
        in_img_array[16][3] <= 18'd0;\
        in_img_array[16][4] <= 18'd0;\
        in_img_array[16][5] <= 18'd0;\
        in_img_array[16][6] <= 18'd0;\
        in_img_array[16][7] <= 18'd0;\
        in_img_array[16][8] <= 18'd0;\
        in_img_array[16][9] <= 18'd0;\
        in_img_array[16][10] <= 18'd0;\
        in_img_array[16][11] <= 18'd0;\
        in_img_array[16][12] <= 18'd0;\
        in_img_array[16][13] <= 18'd0;\
        in_img_array[16][14] <= 18'd0;\
        in_img_array[16][15] <= 18'd0;\
        in_img_array[16][16] <= 18'd0;\
        in_img_array[16][17] <= 18'd0;\
        in_img_array[16][18] <= 18'd0;\
        in_img_array[16][19] <= 18'd0;\
        in_img_array[16][20] <= 18'd0;\
        in_img_array[16][21] <= 18'd0;\
        in_img_array[16][22] <= 18'd0;\
        in_img_array[16][23] <= 18'd0;\
        in_img_array[16][24] <= 18'd0;\
        in_img_array[16][25] <= 18'd0;\
        in_img_array[16][26] <= 18'd0;\
        in_img_array[16][27] <= 18'd0;\
        in_img_array[16][28] <= 18'd0;\
        in_img_array[16][29] <= 18'd0;\
        in_img_array[16][30] <= 18'd0;\
        in_img_array[16][31] <= 18'd0;\
        in_img_array[17][0] <= 18'd0;\
        in_img_array[17][1] <= 18'd0;\
        in_img_array[17][2] <= 18'd0;\
        in_img_array[17][3] <= 18'd0;\
        in_img_array[17][4] <= 18'd0;\
        in_img_array[17][5] <= 18'd0;\
        in_img_array[17][6] <= 18'd0;\
        in_img_array[17][7] <= 18'd0;\
        in_img_array[17][8] <= 18'd0;\
        in_img_array[17][9] <= 18'd0;\
        in_img_array[17][10] <= 18'd0;\
        in_img_array[17][11] <= 18'd0;\
        in_img_array[17][12] <= 18'd0;\
        in_img_array[17][13] <= 18'd0;\
        in_img_array[17][14] <= 18'd0;\
        in_img_array[17][15] <= 18'd0;\
        in_img_array[17][16] <= 18'd0;\
        in_img_array[17][17] <= 18'd0;\
        in_img_array[17][18] <= 18'd0;\
        in_img_array[17][19] <= 18'd0;\
        in_img_array[17][20] <= 18'd0;\
        in_img_array[17][21] <= 18'd0;\
        in_img_array[17][22] <= 18'd0;\
        in_img_array[17][23] <= 18'd0;\
        in_img_array[17][24] <= 18'd0;\
        in_img_array[17][25] <= 18'd0;\
        in_img_array[17][26] <= 18'd0;\
        in_img_array[17][27] <= 18'd0;\
        in_img_array[17][28] <= 18'd0;\
        in_img_array[17][29] <= 18'd0;\
        in_img_array[17][30] <= 18'd0;\
        in_img_array[17][31] <= 18'd0;\
        in_img_array[18][0] <= 18'd0;\
        in_img_array[18][1] <= 18'd0;\
        in_img_array[18][2] <= 18'd0;\
        in_img_array[18][3] <= 18'd0;\
        in_img_array[18][4] <= 18'd0;\
        in_img_array[18][5] <= 18'd0;\
        in_img_array[18][6] <= 18'd0;\
        in_img_array[18][7] <= 18'd0;\
        in_img_array[18][8] <= 18'd0;\
        in_img_array[18][9] <= 18'd0;\
        in_img_array[18][10] <= 18'd0;\
        in_img_array[18][11] <= 18'd0;\
        in_img_array[18][12] <= 18'd0;\
        in_img_array[18][13] <= 18'd0;\
        in_img_array[18][14] <= 18'd0;\
        in_img_array[18][15] <= 18'd0;\
        in_img_array[18][16] <= 18'd0;\
        in_img_array[18][17] <= 18'd0;\
        in_img_array[18][18] <= 18'd0;\
        in_img_array[18][19] <= 18'd0;\
        in_img_array[18][20] <= 18'd0;\
        in_img_array[18][21] <= 18'd0;\
        in_img_array[18][22] <= 18'd0;\
        in_img_array[18][23] <= 18'd0;\
        in_img_array[18][24] <= 18'd0;\
        in_img_array[18][25] <= 18'd0;\
        in_img_array[18][26] <= 18'd0;\
        in_img_array[18][27] <= 18'd0;\
        in_img_array[18][28] <= 18'd0;\
        in_img_array[18][29] <= 18'd0;\
        in_img_array[18][30] <= 18'd0;\
        in_img_array[18][31] <= 18'd0;\
        in_img_array[19][0] <= 18'd0;\
        in_img_array[19][1] <= 18'd0;\
        in_img_array[19][2] <= 18'd0;\
        in_img_array[19][3] <= 18'd0;\
        in_img_array[19][4] <= 18'd0;\
        in_img_array[19][5] <= 18'd0;\
        in_img_array[19][6] <= 18'd0;\
        in_img_array[19][7] <= 18'd0;\
        in_img_array[19][8] <= 18'd0;\
        in_img_array[19][9] <= 18'd0;\
        in_img_array[19][10] <= 18'd0;\
        in_img_array[19][11] <= 18'd0;\
        in_img_array[19][12] <= 18'd0;\
        in_img_array[19][13] <= 18'd0;\
        in_img_array[19][14] <= 18'd0;\
        in_img_array[19][15] <= 18'd0;\
        in_img_array[19][16] <= 18'd0;\
        in_img_array[19][17] <= 18'd0;\
        in_img_array[19][18] <= 18'd0;\
        in_img_array[19][19] <= 18'd0;\
        in_img_array[19][20] <= 18'd0;\
        in_img_array[19][21] <= 18'd0;\
        in_img_array[19][22] <= 18'd0;\
        in_img_array[19][23] <= 18'd0;\
        in_img_array[19][24] <= 18'd0;\
        in_img_array[19][25] <= 18'd0;\
        in_img_array[19][26] <= 18'd0;\
        in_img_array[19][27] <= 18'd0;\
        in_img_array[19][28] <= 18'd0;\
        in_img_array[19][29] <= 18'd0;\
        in_img_array[19][30] <= 18'd0;\
        in_img_array[19][31] <= 18'd0;\
        in_img_array[20][0] <= 18'd0;\
        in_img_array[20][1] <= 18'd0;\
        in_img_array[20][2] <= 18'd0;\
        in_img_array[20][3] <= 18'd0;\
        in_img_array[20][4] <= 18'd0;\
        in_img_array[20][5] <= 18'd0;\
        in_img_array[20][6] <= 18'd0;\
        in_img_array[20][7] <= 18'd0;\
        in_img_array[20][8] <= 18'd0;\
        in_img_array[20][9] <= 18'd0;\
        in_img_array[20][10] <= 18'd0;\
        in_img_array[20][11] <= 18'd0;\
        in_img_array[20][12] <= 18'd0;\
        in_img_array[20][13] <= 18'd0;\
        in_img_array[20][14] <= 18'd0;\
        in_img_array[20][15] <= 18'd0;\
        in_img_array[20][16] <= 18'd0;\
        in_img_array[20][17] <= 18'd0;\
        in_img_array[20][18] <= 18'd0;\
        in_img_array[20][19] <= 18'd0;\
        in_img_array[20][20] <= 18'd0;\
        in_img_array[20][21] <= 18'd0;\
        in_img_array[20][22] <= 18'd0;\
        in_img_array[20][23] <= 18'd0;\
        in_img_array[20][24] <= 18'd0;\
        in_img_array[20][25] <= 18'd0;\
        in_img_array[20][26] <= 18'd0;\
        in_img_array[20][27] <= 18'd0;\
        in_img_array[20][28] <= 18'd0;\
        in_img_array[20][29] <= 18'd0;\
        in_img_array[20][30] <= 18'd0;\
        in_img_array[20][31] <= 18'd0;\
        in_img_array[21][0] <= 18'd0;\
        in_img_array[21][1] <= 18'd0;\
        in_img_array[21][2] <= 18'd0;\
        in_img_array[21][3] <= 18'd0;\
        in_img_array[21][4] <= 18'd0;\
        in_img_array[21][5] <= 18'd0;\
        in_img_array[21][6] <= 18'd0;\
        in_img_array[21][7] <= 18'd0;\
        in_img_array[21][8] <= 18'd0;\
        in_img_array[21][9] <= 18'd0;\
        in_img_array[21][10] <= 18'd0;\
        in_img_array[21][11] <= 18'd0;\
        in_img_array[21][12] <= 18'd0;\
        in_img_array[21][13] <= 18'd0;\
        in_img_array[21][14] <= 18'd0;\
        in_img_array[21][15] <= 18'd0;\
        in_img_array[21][16] <= 18'd0;\
        in_img_array[21][17] <= 18'd0;\
        in_img_array[21][18] <= 18'd0;\
        in_img_array[21][19] <= 18'd0;\
        in_img_array[21][20] <= 18'd0;\
        in_img_array[21][21] <= 18'd0;\
        in_img_array[21][22] <= 18'd0;\
        in_img_array[21][23] <= 18'd0;\
        in_img_array[21][24] <= 18'd0;\
        in_img_array[21][25] <= 18'd0;\
        in_img_array[21][26] <= 18'd0;\
        in_img_array[21][27] <= 18'd0;\
        in_img_array[21][28] <= 18'd0;\
        in_img_array[21][29] <= 18'd0;\
        in_img_array[21][30] <= 18'd0;\
        in_img_array[21][31] <= 18'd0;\
        in_img_array[22][0] <= 18'd0;\
        in_img_array[22][1] <= 18'd0;\
        in_img_array[22][2] <= 18'd0;\
        in_img_array[22][3] <= 18'd0;\
        in_img_array[22][4] <= 18'd0;\
        in_img_array[22][5] <= 18'd0;\
        in_img_array[22][6] <= 18'd0;\
        in_img_array[22][7] <= 18'd0;\
        in_img_array[22][8] <= 18'd0;\
        in_img_array[22][9] <= 18'd0;\
        in_img_array[22][10] <= 18'd0;\
        in_img_array[22][11] <= 18'd0;\
        in_img_array[22][12] <= 18'd0;\
        in_img_array[22][13] <= 18'd0;\
        in_img_array[22][14] <= 18'd0;\
        in_img_array[22][15] <= 18'd0;\
        in_img_array[22][16] <= 18'd0;\
        in_img_array[22][17] <= 18'd0;\
        in_img_array[22][18] <= 18'd0;\
        in_img_array[22][19] <= 18'd0;\
        in_img_array[22][20] <= 18'd0;\
        in_img_array[22][21] <= 18'd0;\
        in_img_array[22][22] <= 18'd0;\
        in_img_array[22][23] <= 18'd0;\
        in_img_array[22][24] <= 18'd0;\
        in_img_array[22][25] <= 18'd0;\
        in_img_array[22][26] <= 18'd0;\
        in_img_array[22][27] <= 18'd0;\
        in_img_array[22][28] <= 18'd0;\
        in_img_array[22][29] <= 18'd0;\
        in_img_array[22][30] <= 18'd0;\
        in_img_array[22][31] <= 18'd0;\
        in_img_array[23][0] <= 18'd0;\
        in_img_array[23][1] <= 18'd0;\
        in_img_array[23][2] <= 18'd0;\
        in_img_array[23][3] <= 18'd0;\
        in_img_array[23][4] <= 18'd0;\
        in_img_array[23][5] <= 18'd0;\
        in_img_array[23][6] <= 18'd0;\
        in_img_array[23][7] <= 18'd0;\
        in_img_array[23][8] <= 18'd0;\
        in_img_array[23][9] <= 18'd0;\
        in_img_array[23][10] <= 18'd0;\
        in_img_array[23][11] <= 18'd0;\
        in_img_array[23][12] <= 18'd0;\
        in_img_array[23][13] <= 18'd0;\
        in_img_array[23][14] <= 18'd0;\
        in_img_array[23][15] <= 18'd0;\
        in_img_array[23][16] <= 18'd0;\
        in_img_array[23][17] <= 18'd0;\
        in_img_array[23][18] <= 18'd0;\
        in_img_array[23][19] <= 18'd0;\
        in_img_array[23][20] <= 18'd0;\
        in_img_array[23][21] <= 18'd0;\
        in_img_array[23][22] <= 18'd0;\
        in_img_array[23][23] <= 18'd0;\
        in_img_array[23][24] <= 18'd0;\
        in_img_array[23][25] <= 18'd0;\
        in_img_array[23][26] <= 18'd0;\
        in_img_array[23][27] <= 18'd0;\
        in_img_array[23][28] <= 18'd0;\
        in_img_array[23][29] <= 18'd0;\
        in_img_array[23][30] <= 18'd0;\
        in_img_array[23][31] <= 18'd0;\
        in_img_array[24][0] <= 18'd0;\
        in_img_array[24][1] <= 18'd0;\
        in_img_array[24][2] <= 18'd0;\
        in_img_array[24][3] <= 18'd0;\
        in_img_array[24][4] <= 18'd0;\
        in_img_array[24][5] <= 18'd0;\
        in_img_array[24][6] <= 18'd0;\
        in_img_array[24][7] <= 18'd0;\
        in_img_array[24][8] <= 18'd0;\
        in_img_array[24][9] <= 18'd0;\
        in_img_array[24][10] <= 18'd0;\
        in_img_array[24][11] <= 18'd0;\
        in_img_array[24][12] <= 18'd0;\
        in_img_array[24][13] <= 18'd0;\
        in_img_array[24][14] <= 18'd0;\
        in_img_array[24][15] <= 18'd0;\
        in_img_array[24][16] <= 18'd0;\
        in_img_array[24][17] <= 18'd0;\
        in_img_array[24][18] <= 18'd0;\
        in_img_array[24][19] <= 18'd0;\
        in_img_array[24][20] <= 18'd0;\
        in_img_array[24][21] <= 18'd0;\
        in_img_array[24][22] <= 18'd0;\
        in_img_array[24][23] <= 18'd0;\
        in_img_array[24][24] <= 18'd0;\
        in_img_array[24][25] <= 18'd0;\
        in_img_array[24][26] <= 18'd0;\
        in_img_array[24][27] <= 18'd0;\
        in_img_array[24][28] <= 18'd0;\
        in_img_array[24][29] <= 18'd0;\
        in_img_array[24][30] <= 18'd0;\
        in_img_array[24][31] <= 18'd0;\
        in_img_array[25][0] <= 18'd0;\
        in_img_array[25][1] <= 18'd0;\
        in_img_array[25][2] <= 18'd0;\
        in_img_array[25][3] <= 18'd0;\
        in_img_array[25][4] <= 18'd0;\
        in_img_array[25][5] <= 18'd0;\
        in_img_array[25][6] <= 18'd0;\
        in_img_array[25][7] <= 18'd0;\
        in_img_array[25][8] <= 18'd0;\
        in_img_array[25][9] <= 18'd0;\
        in_img_array[25][10] <= 18'd0;\
        in_img_array[25][11] <= 18'd0;\
        in_img_array[25][12] <= 18'd0;\
        in_img_array[25][13] <= 18'd0;\
        in_img_array[25][14] <= 18'd0;\
        in_img_array[25][15] <= 18'd0;\
        in_img_array[25][16] <= 18'd0;\
        in_img_array[25][17] <= 18'd0;\
        in_img_array[25][18] <= 18'd0;\
        in_img_array[25][19] <= 18'd0;\
        in_img_array[25][20] <= 18'd0;\
        in_img_array[25][21] <= 18'd0;\
        in_img_array[25][22] <= 18'd0;\
        in_img_array[25][23] <= 18'd0;\
        in_img_array[25][24] <= 18'd0;\
        in_img_array[25][25] <= 18'd0;\
        in_img_array[25][26] <= 18'd0;\
        in_img_array[25][27] <= 18'd0;\
        in_img_array[25][28] <= 18'd0;\
        in_img_array[25][29] <= 18'd0;\
        in_img_array[25][30] <= 18'd0;\
        in_img_array[25][31] <= 18'd0;\
        in_img_array[26][0] <= 18'd0;\
        in_img_array[26][1] <= 18'd0;\
        in_img_array[26][2] <= 18'd0;\
        in_img_array[26][3] <= 18'd0;\
        in_img_array[26][4] <= 18'd0;\
        in_img_array[26][5] <= 18'd0;\
        in_img_array[26][6] <= 18'd0;\
        in_img_array[26][7] <= 18'd0;\
        in_img_array[26][8] <= 18'd0;\
        in_img_array[26][9] <= 18'd0;\
        in_img_array[26][10] <= 18'd0;\
        in_img_array[26][11] <= 18'd0;\
        in_img_array[26][12] <= 18'd0;\
        in_img_array[26][13] <= 18'd0;\
        in_img_array[26][14] <= 18'd0;\
        in_img_array[26][15] <= 18'd0;\
        in_img_array[26][16] <= 18'd0;\
        in_img_array[26][17] <= 18'd0;\
        in_img_array[26][18] <= 18'd0;\
        in_img_array[26][19] <= 18'd0;\
        in_img_array[26][20] <= 18'd0;\
        in_img_array[26][21] <= 18'd0;\
        in_img_array[26][22] <= 18'd0;\
        in_img_array[26][23] <= 18'd0;\
        in_img_array[26][24] <= 18'd0;\
        in_img_array[26][25] <= 18'd0;\
        in_img_array[26][26] <= 18'd0;\
        in_img_array[26][27] <= 18'd0;\
        in_img_array[26][28] <= 18'd0;\
        in_img_array[26][29] <= 18'd0;\
        in_img_array[26][30] <= 18'd0;\
        in_img_array[26][31] <= 18'd0;\
        in_img_array[27][0] <= 18'd0;\
        in_img_array[27][1] <= 18'd0;\
        in_img_array[27][2] <= 18'd0;\
        in_img_array[27][3] <= 18'd0;\
        in_img_array[27][4] <= 18'd0;\
        in_img_array[27][5] <= 18'd0;\
        in_img_array[27][6] <= 18'd0;\
        in_img_array[27][7] <= 18'd0;\
        in_img_array[27][8] <= 18'd0;\
        in_img_array[27][9] <= 18'd0;\
        in_img_array[27][10] <= 18'd0;\
        in_img_array[27][11] <= 18'd0;\
        in_img_array[27][12] <= 18'd0;\
        in_img_array[27][13] <= 18'd0;\
        in_img_array[27][14] <= 18'd0;\
        in_img_array[27][15] <= 18'd0;\
        in_img_array[27][16] <= 18'd0;\
        in_img_array[27][17] <= 18'd0;\
        in_img_array[27][18] <= 18'd0;\
        in_img_array[27][19] <= 18'd0;\
        in_img_array[27][20] <= 18'd0;\
        in_img_array[27][21] <= 18'd0;\
        in_img_array[27][22] <= 18'd0;\
        in_img_array[27][23] <= 18'd0;\
        in_img_array[27][24] <= 18'd0;\
        in_img_array[27][25] <= 18'd0;\
        in_img_array[27][26] <= 18'd0;\
        in_img_array[27][27] <= 18'd0;\
        in_img_array[27][28] <= 18'd0;\
        in_img_array[27][29] <= 18'd0;\
        in_img_array[27][30] <= 18'd0;\
        in_img_array[27][31] <= 18'd0;\
        in_img_array[28][0] <= 18'd0;\
        in_img_array[28][1] <= 18'd0;\
        in_img_array[28][2] <= 18'd0;\
        in_img_array[28][3] <= 18'd0;\
        in_img_array[28][4] <= 18'd0;\
        in_img_array[28][5] <= 18'd0;\
        in_img_array[28][6] <= 18'd0;\
        in_img_array[28][7] <= 18'd0;\
        in_img_array[28][8] <= 18'd0;\
        in_img_array[28][9] <= 18'd0;\
        in_img_array[28][10] <= 18'd0;\
        in_img_array[28][11] <= 18'd0;\
        in_img_array[28][12] <= 18'd0;\
        in_img_array[28][13] <= 18'd0;\
        in_img_array[28][14] <= 18'd0;\
        in_img_array[28][15] <= 18'd0;\
        in_img_array[28][16] <= 18'd0;\
        in_img_array[28][17] <= 18'd0;\
        in_img_array[28][18] <= 18'd0;\
        in_img_array[28][19] <= 18'd0;\
        in_img_array[28][20] <= 18'd0;\
        in_img_array[28][21] <= 18'd0;\
        in_img_array[28][22] <= 18'd0;\
        in_img_array[28][23] <= 18'd0;\
        in_img_array[28][24] <= 18'd0;\
        in_img_array[28][25] <= 18'd0;\
        in_img_array[28][26] <= 18'd0;\
        in_img_array[28][27] <= 18'd0;\
        in_img_array[28][28] <= 18'd0;\
        in_img_array[28][29] <= 18'd0;\
        in_img_array[28][30] <= 18'd0;\
        in_img_array[28][31] <= 18'd0;\
        in_img_array[29][0] <= 18'd0;\
        in_img_array[29][1] <= 18'd0;\
        in_img_array[29][2] <= 18'd0;\
        in_img_array[29][3] <= 18'd0;\
        in_img_array[29][4] <= 18'd0;\
        in_img_array[29][5] <= 18'd0;\
        in_img_array[29][6] <= 18'd0;\
        in_img_array[29][7] <= 18'd0;\
        in_img_array[29][8] <= 18'd0;\
        in_img_array[29][9] <= 18'd0;\
        in_img_array[29][10] <= 18'd0;\
        in_img_array[29][11] <= 18'd0;\
        in_img_array[29][12] <= 18'd0;\
        in_img_array[29][13] <= 18'd0;\
        in_img_array[29][14] <= 18'd0;\
        in_img_array[29][15] <= 18'd0;\
        in_img_array[29][16] <= 18'd0;\
        in_img_array[29][17] <= 18'd0;\
        in_img_array[29][18] <= 18'd0;\
        in_img_array[29][19] <= 18'd0;\
        in_img_array[29][20] <= 18'd0;\
        in_img_array[29][21] <= 18'd0;\
        in_img_array[29][22] <= 18'd0;\
        in_img_array[29][23] <= 18'd0;\
        in_img_array[29][24] <= 18'd0;\
        in_img_array[29][25] <= 18'd0;\
        in_img_array[29][26] <= 18'd0;\
        in_img_array[29][27] <= 18'd0;\
        in_img_array[29][28] <= 18'd0;\
        in_img_array[29][29] <= 18'd0;\
        in_img_array[29][30] <= 18'd0;\
        in_img_array[29][31] <= 18'd0;\
        in_img_array[30][0] <= 18'd0;\
        in_img_array[30][1] <= 18'd0;\
        in_img_array[30][2] <= 18'd0;\
        in_img_array[30][3] <= 18'd0;\
        in_img_array[30][4] <= 18'd0;\
        in_img_array[30][5] <= 18'd0;\
        in_img_array[30][6] <= 18'd0;\
        in_img_array[30][7] <= 18'd0;\
        in_img_array[30][8] <= 18'd0;\
        in_img_array[30][9] <= 18'd0;\
        in_img_array[30][10] <= 18'd0;\
        in_img_array[30][11] <= 18'd0;\
        in_img_array[30][12] <= 18'd0;\
        in_img_array[30][13] <= 18'd0;\
        in_img_array[30][14] <= 18'd0;\
        in_img_array[30][15] <= 18'd0;\
        in_img_array[30][16] <= 18'd0;\
        in_img_array[30][17] <= 18'd0;\
        in_img_array[30][18] <= 18'd0;\
        in_img_array[30][19] <= 18'd0;\
        in_img_array[30][20] <= 18'd0;\
        in_img_array[30][21] <= 18'd0;\
        in_img_array[30][22] <= 18'd0;\
        in_img_array[30][23] <= 18'd0;\
        in_img_array[30][24] <= 18'd0;\
        in_img_array[30][25] <= 18'd0;\
        in_img_array[30][26] <= 18'd0;\
        in_img_array[30][27] <= 18'd0;\
        in_img_array[30][28] <= 18'd0;\
        in_img_array[30][29] <= 18'd0;\
        in_img_array[30][30] <= 18'd0;\
        in_img_array[30][31] <= 18'd0;\
        in_img_array[31][0] <= 18'd0;\
        in_img_array[31][1] <= 18'd0;\
        in_img_array[31][2] <= 18'd0;\
        in_img_array[31][3] <= 18'd0;\
        in_img_array[31][4] <= 18'd0;\
        in_img_array[31][5] <= 18'd0;\
        in_img_array[31][6] <= 18'd0;\
        in_img_array[31][7] <= 18'd0;\
        in_img_array[31][8] <= 18'd0;\
        in_img_array[31][9] <= 18'd0;\
        in_img_array[31][10] <= 18'd0;\
        in_img_array[31][11] <= 18'd0;\
        in_img_array[31][12] <= 18'd0;\
        in_img_array[31][13] <= 18'd0;\
        in_img_array[31][14] <= 18'd0;\
        in_img_array[31][15] <= 18'd0;\
        in_img_array[31][16] <= 18'd0;\
        in_img_array[31][17] <= 18'd0;\
        in_img_array[31][18] <= 18'd0;\
        in_img_array[31][19] <= 18'd0;\
        in_img_array[31][20] <= 18'd0;\
        in_img_array[31][21] <= 18'd0;\
        in_img_array[31][22] <= 18'd0;\
        in_img_array[31][23] <= 18'd0;\
        in_img_array[31][24] <= 18'd0;\
        in_img_array[31][25] <= 18'd0;\
        in_img_array[31][26] <= 18'd0;\
        in_img_array[31][27] <= 18'd0;\
        in_img_array[31][28] <= 18'd0;\
        in_img_array[31][29] <= 18'd0;\
        in_img_array[31][30] <= 18'd0;\
        in_img_array[31][31] <= 18'd0;\
    end\
    else if((state==IDLE)&(pre_finish))begin\
        in_img_array[2][2][0] <= img[0];\
        in_img_array[2][2][1] <= img[1];\
        in_img_array[2][2][2] <= img[2];\
        in_img_array[2][2][3] <= img[3];\
        in_img_array[2][2][4] <= img[4];\
        in_img_array[2][2][5] <= img[5];\
        in_img_array[2][2][6] <= img[6];\
        in_img_array[2][2][7] <= img[7];\
        in_img_array[2][2][8] <= img[8];\
        in_img_array[2][2][9] <= img[9];\
        in_img_array[2][2][10] <= img[10];\
        in_img_array[2][2][11] <= img[11];\
        in_img_array[2][2][12] <= img[12];\
        in_img_array[2][2][13] <= img[13];\
        in_img_array[2][2][14] <= img[14];\
        in_img_array[2][2][15] <= img[15];\
        in_img_array[2][2][16] <= img[16];\
        in_img_array[2][2][17] <= img[17];\
        in_img_array[2][3][0] <= img[18];\
        in_img_array[2][3][1] <= img[19];\
        in_img_array[2][3][2] <= img[20];\
        in_img_array[2][3][3] <= img[21];\
        in_img_array[2][3][4] <= img[22];\
        in_img_array[2][3][5] <= img[23];\
        in_img_array[2][3][6] <= img[24];\
        in_img_array[2][3][7] <= img[25];\
        in_img_array[2][3][8] <= img[26];\
        in_img_array[2][3][9] <= img[27];\
        in_img_array[2][3][10] <= img[28];\
        in_img_array[2][3][11] <= img[29];\
        in_img_array[2][3][12] <= img[30];\
        in_img_array[2][3][13] <= img[31];\
        in_img_array[2][3][14] <= img[32];\
        in_img_array[2][3][15] <= img[33];\
        in_img_array[2][3][16] <= img[34];\
        in_img_array[2][3][17] <= img[35];\
        in_img_array[2][4][0] <= img[36];\
        in_img_array[2][4][1] <= img[37];\
        in_img_array[2][4][2] <= img[38];\
        in_img_array[2][4][3] <= img[39];\
        in_img_array[2][4][4] <= img[40];\
        in_img_array[2][4][5] <= img[41];\
        in_img_array[2][4][6] <= img[42];\
        in_img_array[2][4][7] <= img[43];\
        in_img_array[2][4][8] <= img[44];\
        in_img_array[2][4][9] <= img[45];\
        in_img_array[2][4][10] <= img[46];\
        in_img_array[2][4][11] <= img[47];\
        in_img_array[2][4][12] <= img[48];\
        in_img_array[2][4][13] <= img[49];\
        in_img_array[2][4][14] <= img[50];\
        in_img_array[2][4][15] <= img[51];\
        in_img_array[2][4][16] <= img[52];\
        in_img_array[2][4][17] <= img[53];\
        in_img_array[2][5][0] <= img[54];\
        in_img_array[2][5][1] <= img[55];\
        in_img_array[2][5][2] <= img[56];\
        in_img_array[2][5][3] <= img[57];\
        in_img_array[2][5][4] <= img[58];\
        in_img_array[2][5][5] <= img[59];\
        in_img_array[2][5][6] <= img[60];\
        in_img_array[2][5][7] <= img[61];\
        in_img_array[2][5][8] <= img[62];\
        in_img_array[2][5][9] <= img[63];\
        in_img_array[2][5][10] <= img[64];\
        in_img_array[2][5][11] <= img[65];\
        in_img_array[2][5][12] <= img[66];\
        in_img_array[2][5][13] <= img[67];\
        in_img_array[2][5][14] <= img[68];\
        in_img_array[2][5][15] <= img[69];\
        in_img_array[2][5][16] <= img[70];\
        in_img_array[2][5][17] <= img[71];\
        in_img_array[2][6][0] <= img[72];\
        in_img_array[2][6][1] <= img[73];\
        in_img_array[2][6][2] <= img[74];\
        in_img_array[2][6][3] <= img[75];\
        in_img_array[2][6][4] <= img[76];\
        in_img_array[2][6][5] <= img[77];\
        in_img_array[2][6][6] <= img[78];\
        in_img_array[2][6][7] <= img[79];\
        in_img_array[2][6][8] <= img[80];\
        in_img_array[2][6][9] <= img[81];\
        in_img_array[2][6][10] <= img[82];\
        in_img_array[2][6][11] <= img[83];\
        in_img_array[2][6][12] <= img[84];\
        in_img_array[2][6][13] <= img[85];\
        in_img_array[2][6][14] <= img[86];\
        in_img_array[2][6][15] <= img[87];\
        in_img_array[2][6][16] <= img[88];\
        in_img_array[2][6][17] <= img[89];\
        in_img_array[2][7][0] <= img[90];\
        in_img_array[2][7][1] <= img[91];\
        in_img_array[2][7][2] <= img[92];\
        in_img_array[2][7][3] <= img[93];\
        in_img_array[2][7][4] <= img[94];\
        in_img_array[2][7][5] <= img[95];\
        in_img_array[2][7][6] <= img[96];\
        in_img_array[2][7][7] <= img[97];\
        in_img_array[2][7][8] <= img[98];\
        in_img_array[2][7][9] <= img[99];\
        in_img_array[2][7][10] <= img[100];\
        in_img_array[2][7][11] <= img[101];\
        in_img_array[2][7][12] <= img[102];\
        in_img_array[2][7][13] <= img[103];\
        in_img_array[2][7][14] <= img[104];\
        in_img_array[2][7][15] <= img[105];\
        in_img_array[2][7][16] <= img[106];\
        in_img_array[2][7][17] <= img[107];\
        in_img_array[2][8][0] <= img[108];\
        in_img_array[2][8][1] <= img[109];\
        in_img_array[2][8][2] <= img[110];\
        in_img_array[2][8][3] <= img[111];\
        in_img_array[2][8][4] <= img[112];\
        in_img_array[2][8][5] <= img[113];\
        in_img_array[2][8][6] <= img[114];\
        in_img_array[2][8][7] <= img[115];\
        in_img_array[2][8][8] <= img[116];\
        in_img_array[2][8][9] <= img[117];\
        in_img_array[2][8][10] <= img[118];\
        in_img_array[2][8][11] <= img[119];\
        in_img_array[2][8][12] <= img[120];\
        in_img_array[2][8][13] <= img[121];\
        in_img_array[2][8][14] <= img[122];\
        in_img_array[2][8][15] <= img[123];\
        in_img_array[2][8][16] <= img[124];\
        in_img_array[2][8][17] <= img[125];\
        in_img_array[2][9][0] <= img[126];\
        in_img_array[2][9][1] <= img[127];\
        in_img_array[2][9][2] <= img[128];\
        in_img_array[2][9][3] <= img[129];\
        in_img_array[2][9][4] <= img[130];\
        in_img_array[2][9][5] <= img[131];\
        in_img_array[2][9][6] <= img[132];\
        in_img_array[2][9][7] <= img[133];\
        in_img_array[2][9][8] <= img[134];\
        in_img_array[2][9][9] <= img[135];\
        in_img_array[2][9][10] <= img[136];\
        in_img_array[2][9][11] <= img[137];\
        in_img_array[2][9][12] <= img[138];\
        in_img_array[2][9][13] <= img[139];\
        in_img_array[2][9][14] <= img[140];\
        in_img_array[2][9][15] <= img[141];\
        in_img_array[2][9][16] <= img[142];\
        in_img_array[2][9][17] <= img[143];\
        in_img_array[2][10][0] <= img[144];\
        in_img_array[2][10][1] <= img[145];\
        in_img_array[2][10][2] <= img[146];\
        in_img_array[2][10][3] <= img[147];\
        in_img_array[2][10][4] <= img[148];\
        in_img_array[2][10][5] <= img[149];\
        in_img_array[2][10][6] <= img[150];\
        in_img_array[2][10][7] <= img[151];\
        in_img_array[2][10][8] <= img[152];\
        in_img_array[2][10][9] <= img[153];\
        in_img_array[2][10][10] <= img[154];\
        in_img_array[2][10][11] <= img[155];\
        in_img_array[2][10][12] <= img[156];\
        in_img_array[2][10][13] <= img[157];\
        in_img_array[2][10][14] <= img[158];\
        in_img_array[2][10][15] <= img[159];\
        in_img_array[2][10][16] <= img[160];\
        in_img_array[2][10][17] <= img[161];\
        in_img_array[2][11][0] <= img[162];\
        in_img_array[2][11][1] <= img[163];\
        in_img_array[2][11][2] <= img[164];\
        in_img_array[2][11][3] <= img[165];\
        in_img_array[2][11][4] <= img[166];\
        in_img_array[2][11][5] <= img[167];\
        in_img_array[2][11][6] <= img[168];\
        in_img_array[2][11][7] <= img[169];\
        in_img_array[2][11][8] <= img[170];\
        in_img_array[2][11][9] <= img[171];\
        in_img_array[2][11][10] <= img[172];\
        in_img_array[2][11][11] <= img[173];\
        in_img_array[2][11][12] <= img[174];\
        in_img_array[2][11][13] <= img[175];\
        in_img_array[2][11][14] <= img[176];\
        in_img_array[2][11][15] <= img[177];\
        in_img_array[2][11][16] <= img[178];\
        in_img_array[2][11][17] <= img[179];\
        in_img_array[2][12][0] <= img[180];\
        in_img_array[2][12][1] <= img[181];\
        in_img_array[2][12][2] <= img[182];\
        in_img_array[2][12][3] <= img[183];\
        in_img_array[2][12][4] <= img[184];\
        in_img_array[2][12][5] <= img[185];\
        in_img_array[2][12][6] <= img[186];\
        in_img_array[2][12][7] <= img[187];\
        in_img_array[2][12][8] <= img[188];\
        in_img_array[2][12][9] <= img[189];\
        in_img_array[2][12][10] <= img[190];\
        in_img_array[2][12][11] <= img[191];\
        in_img_array[2][12][12] <= img[192];\
        in_img_array[2][12][13] <= img[193];\
        in_img_array[2][12][14] <= img[194];\
        in_img_array[2][12][15] <= img[195];\
        in_img_array[2][12][16] <= img[196];\
        in_img_array[2][12][17] <= img[197];\
        in_img_array[2][13][0] <= img[198];\
        in_img_array[2][13][1] <= img[199];\
        in_img_array[2][13][2] <= img[200];\
        in_img_array[2][13][3] <= img[201];\
        in_img_array[2][13][4] <= img[202];\
        in_img_array[2][13][5] <= img[203];\
        in_img_array[2][13][6] <= img[204];\
        in_img_array[2][13][7] <= img[205];\
        in_img_array[2][13][8] <= img[206];\
        in_img_array[2][13][9] <= img[207];\
        in_img_array[2][13][10] <= img[208];\
        in_img_array[2][13][11] <= img[209];\
        in_img_array[2][13][12] <= img[210];\
        in_img_array[2][13][13] <= img[211];\
        in_img_array[2][13][14] <= img[212];\
        in_img_array[2][13][15] <= img[213];\
        in_img_array[2][13][16] <= img[214];\
        in_img_array[2][13][17] <= img[215];\
        in_img_array[2][14][0] <= img[216];\
        in_img_array[2][14][1] <= img[217];\
        in_img_array[2][14][2] <= img[218];\
        in_img_array[2][14][3] <= img[219];\
        in_img_array[2][14][4] <= img[220];\
        in_img_array[2][14][5] <= img[221];\
        in_img_array[2][14][6] <= img[222];\
        in_img_array[2][14][7] <= img[223];\
        in_img_array[2][14][8] <= img[224];\
        in_img_array[2][14][9] <= img[225];\
        in_img_array[2][14][10] <= img[226];\
        in_img_array[2][14][11] <= img[227];\
        in_img_array[2][14][12] <= img[228];\
        in_img_array[2][14][13] <= img[229];\
        in_img_array[2][14][14] <= img[230];\
        in_img_array[2][14][15] <= img[231];\
        in_img_array[2][14][16] <= img[232];\
        in_img_array[2][14][17] <= img[233];\
        in_img_array[2][15][0] <= img[234];\
        in_img_array[2][15][1] <= img[235];\
        in_img_array[2][15][2] <= img[236];\
        in_img_array[2][15][3] <= img[237];\
        in_img_array[2][15][4] <= img[238];\
        in_img_array[2][15][5] <= img[239];\
        in_img_array[2][15][6] <= img[240];\
        in_img_array[2][15][7] <= img[241];\
        in_img_array[2][15][8] <= img[242];\
        in_img_array[2][15][9] <= img[243];\
        in_img_array[2][15][10] <= img[244];\
        in_img_array[2][15][11] <= img[245];\
        in_img_array[2][15][12] <= img[246];\
        in_img_array[2][15][13] <= img[247];\
        in_img_array[2][15][14] <= img[248];\
        in_img_array[2][15][15] <= img[249];\
        in_img_array[2][15][16] <= img[250];\
        in_img_array[2][15][17] <= img[251];\
        in_img_array[2][16][0] <= img[252];\
        in_img_array[2][16][1] <= img[253];\
        in_img_array[2][16][2] <= img[254];\
        in_img_array[2][16][3] <= img[255];\
        in_img_array[2][16][4] <= img[256];\
        in_img_array[2][16][5] <= img[257];\
        in_img_array[2][16][6] <= img[258];\
        in_img_array[2][16][7] <= img[259];\
        in_img_array[2][16][8] <= img[260];\
        in_img_array[2][16][9] <= img[261];\
        in_img_array[2][16][10] <= img[262];\
        in_img_array[2][16][11] <= img[263];\
        in_img_array[2][16][12] <= img[264];\
        in_img_array[2][16][13] <= img[265];\
        in_img_array[2][16][14] <= img[266];\
        in_img_array[2][16][15] <= img[267];\
        in_img_array[2][16][16] <= img[268];\
        in_img_array[2][16][17] <= img[269];\
        in_img_array[2][17][0] <= img[270];\
        in_img_array[2][17][1] <= img[271];\
        in_img_array[2][17][2] <= img[272];\
        in_img_array[2][17][3] <= img[273];\
        in_img_array[2][17][4] <= img[274];\
        in_img_array[2][17][5] <= img[275];\
        in_img_array[2][17][6] <= img[276];\
        in_img_array[2][17][7] <= img[277];\
        in_img_array[2][17][8] <= img[278];\
        in_img_array[2][17][9] <= img[279];\
        in_img_array[2][17][10] <= img[280];\
        in_img_array[2][17][11] <= img[281];\
        in_img_array[2][17][12] <= img[282];\
        in_img_array[2][17][13] <= img[283];\
        in_img_array[2][17][14] <= img[284];\
        in_img_array[2][17][15] <= img[285];\
        in_img_array[2][17][16] <= img[286];\
        in_img_array[2][17][17] <= img[287];\
        in_img_array[2][18][0] <= img[288];\
        in_img_array[2][18][1] <= img[289];\
        in_img_array[2][18][2] <= img[290];\
        in_img_array[2][18][3] <= img[291];\
        in_img_array[2][18][4] <= img[292];\
        in_img_array[2][18][5] <= img[293];\
        in_img_array[2][18][6] <= img[294];\
        in_img_array[2][18][7] <= img[295];\
        in_img_array[2][18][8] <= img[296];\
        in_img_array[2][18][9] <= img[297];\
        in_img_array[2][18][10] <= img[298];\
        in_img_array[2][18][11] <= img[299];\
        in_img_array[2][18][12] <= img[300];\
        in_img_array[2][18][13] <= img[301];\
        in_img_array[2][18][14] <= img[302];\
        in_img_array[2][18][15] <= img[303];\
        in_img_array[2][18][16] <= img[304];\
        in_img_array[2][18][17] <= img[305];\
        in_img_array[2][19][0] <= img[306];\
        in_img_array[2][19][1] <= img[307];\
        in_img_array[2][19][2] <= img[308];\
        in_img_array[2][19][3] <= img[309];\
        in_img_array[2][19][4] <= img[310];\
        in_img_array[2][19][5] <= img[311];\
        in_img_array[2][19][6] <= img[312];\
        in_img_array[2][19][7] <= img[313];\
        in_img_array[2][19][8] <= img[314];\
        in_img_array[2][19][9] <= img[315];\
        in_img_array[2][19][10] <= img[316];\
        in_img_array[2][19][11] <= img[317];\
        in_img_array[2][19][12] <= img[318];\
        in_img_array[2][19][13] <= img[319];\
        in_img_array[2][19][14] <= img[320];\
        in_img_array[2][19][15] <= img[321];\
        in_img_array[2][19][16] <= img[322];\
        in_img_array[2][19][17] <= img[323];\
        in_img_array[2][20][0] <= img[324];\
        in_img_array[2][20][1] <= img[325];\
        in_img_array[2][20][2] <= img[326];\
        in_img_array[2][20][3] <= img[327];\
        in_img_array[2][20][4] <= img[328];\
        in_img_array[2][20][5] <= img[329];\
        in_img_array[2][20][6] <= img[330];\
        in_img_array[2][20][7] <= img[331];\
        in_img_array[2][20][8] <= img[332];\
        in_img_array[2][20][9] <= img[333];\
        in_img_array[2][20][10] <= img[334];\
        in_img_array[2][20][11] <= img[335];\
        in_img_array[2][20][12] <= img[336];\
        in_img_array[2][20][13] <= img[337];\
        in_img_array[2][20][14] <= img[338];\
        in_img_array[2][20][15] <= img[339];\
        in_img_array[2][20][16] <= img[340];\
        in_img_array[2][20][17] <= img[341];\
        in_img_array[2][21][0] <= img[342];\
        in_img_array[2][21][1] <= img[343];\
        in_img_array[2][21][2] <= img[344];\
        in_img_array[2][21][3] <= img[345];\
        in_img_array[2][21][4] <= img[346];\
        in_img_array[2][21][5] <= img[347];\
        in_img_array[2][21][6] <= img[348];\
        in_img_array[2][21][7] <= img[349];\
        in_img_array[2][21][8] <= img[350];\
        in_img_array[2][21][9] <= img[351];\
        in_img_array[2][21][10] <= img[352];\
        in_img_array[2][21][11] <= img[353];\
        in_img_array[2][21][12] <= img[354];\
        in_img_array[2][21][13] <= img[355];\
        in_img_array[2][21][14] <= img[356];\
        in_img_array[2][21][15] <= img[357];\
        in_img_array[2][21][16] <= img[358];\
        in_img_array[2][21][17] <= img[359];\
        in_img_array[2][22][0] <= img[360];\
        in_img_array[2][22][1] <= img[361];\
        in_img_array[2][22][2] <= img[362];\
        in_img_array[2][22][3] <= img[363];\
        in_img_array[2][22][4] <= img[364];\
        in_img_array[2][22][5] <= img[365];\
        in_img_array[2][22][6] <= img[366];\
        in_img_array[2][22][7] <= img[367];\
        in_img_array[2][22][8] <= img[368];\
        in_img_array[2][22][9] <= img[369];\
        in_img_array[2][22][10] <= img[370];\
        in_img_array[2][22][11] <= img[371];\
        in_img_array[2][22][12] <= img[372];\
        in_img_array[2][22][13] <= img[373];\
        in_img_array[2][22][14] <= img[374];\
        in_img_array[2][22][15] <= img[375];\
        in_img_array[2][22][16] <= img[376];\
        in_img_array[2][22][17] <= img[377];\
        in_img_array[2][23][0] <= img[378];\
        in_img_array[2][23][1] <= img[379];\
        in_img_array[2][23][2] <= img[380];\
        in_img_array[2][23][3] <= img[381];\
        in_img_array[2][23][4] <= img[382];\
        in_img_array[2][23][5] <= img[383];\
        in_img_array[2][23][6] <= img[384];\
        in_img_array[2][23][7] <= img[385];\
        in_img_array[2][23][8] <= img[386];\
        in_img_array[2][23][9] <= img[387];\
        in_img_array[2][23][10] <= img[388];\
        in_img_array[2][23][11] <= img[389];\
        in_img_array[2][23][12] <= img[390];\
        in_img_array[2][23][13] <= img[391];\
        in_img_array[2][23][14] <= img[392];\
        in_img_array[2][23][15] <= img[393];\
        in_img_array[2][23][16] <= img[394];\
        in_img_array[2][23][17] <= img[395];\
        in_img_array[2][24][0] <= img[396];\
        in_img_array[2][24][1] <= img[397];\
        in_img_array[2][24][2] <= img[398];\
        in_img_array[2][24][3] <= img[399];\
        in_img_array[2][24][4] <= img[400];\
        in_img_array[2][24][5] <= img[401];\
        in_img_array[2][24][6] <= img[402];\
        in_img_array[2][24][7] <= img[403];\
        in_img_array[2][24][8] <= img[404];\
        in_img_array[2][24][9] <= img[405];\
        in_img_array[2][24][10] <= img[406];\
        in_img_array[2][24][11] <= img[407];\
        in_img_array[2][24][12] <= img[408];\
        in_img_array[2][24][13] <= img[409];\
        in_img_array[2][24][14] <= img[410];\
        in_img_array[2][24][15] <= img[411];\
        in_img_array[2][24][16] <= img[412];\
        in_img_array[2][24][17] <= img[413];\
        in_img_array[2][25][0] <= img[414];\
        in_img_array[2][25][1] <= img[415];\
        in_img_array[2][25][2] <= img[416];\
        in_img_array[2][25][3] <= img[417];\
        in_img_array[2][25][4] <= img[418];\
        in_img_array[2][25][5] <= img[419];\
        in_img_array[2][25][6] <= img[420];\
        in_img_array[2][25][7] <= img[421];\
        in_img_array[2][25][8] <= img[422];\
        in_img_array[2][25][9] <= img[423];\
        in_img_array[2][25][10] <= img[424];\
        in_img_array[2][25][11] <= img[425];\
        in_img_array[2][25][12] <= img[426];\
        in_img_array[2][25][13] <= img[427];\
        in_img_array[2][25][14] <= img[428];\
        in_img_array[2][25][15] <= img[429];\
        in_img_array[2][25][16] <= img[430];\
        in_img_array[2][25][17] <= img[431];\
        in_img_array[2][26][0] <= img[432];\
        in_img_array[2][26][1] <= img[433];\
        in_img_array[2][26][2] <= img[434];\
        in_img_array[2][26][3] <= img[435];\
        in_img_array[2][26][4] <= img[436];\
        in_img_array[2][26][5] <= img[437];\
        in_img_array[2][26][6] <= img[438];\
        in_img_array[2][26][7] <= img[439];\
        in_img_array[2][26][8] <= img[440];\
        in_img_array[2][26][9] <= img[441];\
        in_img_array[2][26][10] <= img[442];\
        in_img_array[2][26][11] <= img[443];\
        in_img_array[2][26][12] <= img[444];\
        in_img_array[2][26][13] <= img[445];\
        in_img_array[2][26][14] <= img[446];\
        in_img_array[2][26][15] <= img[447];\
        in_img_array[2][26][16] <= img[448];\
        in_img_array[2][26][17] <= img[449];\
        in_img_array[2][27][0] <= img[450];\
        in_img_array[2][27][1] <= img[451];\
        in_img_array[2][27][2] <= img[452];\
        in_img_array[2][27][3] <= img[453];\
        in_img_array[2][27][4] <= img[454];\
        in_img_array[2][27][5] <= img[455];\
        in_img_array[2][27][6] <= img[456];\
        in_img_array[2][27][7] <= img[457];\
        in_img_array[2][27][8] <= img[458];\
        in_img_array[2][27][9] <= img[459];\
        in_img_array[2][27][10] <= img[460];\
        in_img_array[2][27][11] <= img[461];\
        in_img_array[2][27][12] <= img[462];\
        in_img_array[2][27][13] <= img[463];\
        in_img_array[2][27][14] <= img[464];\
        in_img_array[2][27][15] <= img[465];\
        in_img_array[2][27][16] <= img[466];\
        in_img_array[2][27][17] <= img[467];\
        in_img_array[2][28][0] <= img[468];\
        in_img_array[2][28][1] <= img[469];\
        in_img_array[2][28][2] <= img[470];\
        in_img_array[2][28][3] <= img[471];\
        in_img_array[2][28][4] <= img[472];\
        in_img_array[2][28][5] <= img[473];\
        in_img_array[2][28][6] <= img[474];\
        in_img_array[2][28][7] <= img[475];\
        in_img_array[2][28][8] <= img[476];\
        in_img_array[2][28][9] <= img[477];\
        in_img_array[2][28][10] <= img[478];\
        in_img_array[2][28][11] <= img[479];\
        in_img_array[2][28][12] <= img[480];\
        in_img_array[2][28][13] <= img[481];\
        in_img_array[2][28][14] <= img[482];\
        in_img_array[2][28][15] <= img[483];\
        in_img_array[2][28][16] <= img[484];\
        in_img_array[2][28][17] <= img[485];\
        in_img_array[2][29][0] <= img[486];\
        in_img_array[2][29][1] <= img[487];\
        in_img_array[2][29][2] <= img[488];\
        in_img_array[2][29][3] <= img[489];\
        in_img_array[2][29][4] <= img[490];\
        in_img_array[2][29][5] <= img[491];\
        in_img_array[2][29][6] <= img[492];\
        in_img_array[2][29][7] <= img[493];\
        in_img_array[2][29][8] <= img[494];\
        in_img_array[2][29][9] <= img[495];\
        in_img_array[2][29][10] <= img[496];\
        in_img_array[2][29][11] <= img[497];\
        in_img_array[2][29][12] <= img[498];\
        in_img_array[2][29][13] <= img[499];\
        in_img_array[2][29][14] <= img[500];\
        in_img_array[2][29][15] <= img[501];\
        in_img_array[2][29][16] <= img[502];\
        in_img_array[2][29][17] <= img[503];\
        in_img_array[3][2][0] <= img[504];\
        in_img_array[3][2][1] <= img[505];\
        in_img_array[3][2][2] <= img[506];\
        in_img_array[3][2][3] <= img[507];\
        in_img_array[3][2][4] <= img[508];\
        in_img_array[3][2][5] <= img[509];\
        in_img_array[3][2][6] <= img[510];\
        in_img_array[3][2][7] <= img[511];\
        in_img_array[3][2][8] <= img[512];\
        in_img_array[3][2][9] <= img[513];\
        in_img_array[3][2][10] <= img[514];\
        in_img_array[3][2][11] <= img[515];\
        in_img_array[3][2][12] <= img[516];\
        in_img_array[3][2][13] <= img[517];\
        in_img_array[3][2][14] <= img[518];\
        in_img_array[3][2][15] <= img[519];\
        in_img_array[3][2][16] <= img[520];\
        in_img_array[3][2][17] <= img[521];\
        in_img_array[3][3][0] <= img[522];\
        in_img_array[3][3][1] <= img[523];\
        in_img_array[3][3][2] <= img[524];\
        in_img_array[3][3][3] <= img[525];\
        in_img_array[3][3][4] <= img[526];\
        in_img_array[3][3][5] <= img[527];\
        in_img_array[3][3][6] <= img[528];\
        in_img_array[3][3][7] <= img[529];\
        in_img_array[3][3][8] <= img[530];\
        in_img_array[3][3][9] <= img[531];\
        in_img_array[3][3][10] <= img[532];\
        in_img_array[3][3][11] <= img[533];\
        in_img_array[3][3][12] <= img[534];\
        in_img_array[3][3][13] <= img[535];\
        in_img_array[3][3][14] <= img[536];\
        in_img_array[3][3][15] <= img[537];\
        in_img_array[3][3][16] <= img[538];\
        in_img_array[3][3][17] <= img[539];\
        in_img_array[3][4][0] <= img[540];\
        in_img_array[3][4][1] <= img[541];\
        in_img_array[3][4][2] <= img[542];\
        in_img_array[3][4][3] <= img[543];\
        in_img_array[3][4][4] <= img[544];\
        in_img_array[3][4][5] <= img[545];\
        in_img_array[3][4][6] <= img[546];\
        in_img_array[3][4][7] <= img[547];\
        in_img_array[3][4][8] <= img[548];\
        in_img_array[3][4][9] <= img[549];\
        in_img_array[3][4][10] <= img[550];\
        in_img_array[3][4][11] <= img[551];\
        in_img_array[3][4][12] <= img[552];\
        in_img_array[3][4][13] <= img[553];\
        in_img_array[3][4][14] <= img[554];\
        in_img_array[3][4][15] <= img[555];\
        in_img_array[3][4][16] <= img[556];\
        in_img_array[3][4][17] <= img[557];\
        in_img_array[3][5][0] <= img[558];\
        in_img_array[3][5][1] <= img[559];\
        in_img_array[3][5][2] <= img[560];\
        in_img_array[3][5][3] <= img[561];\
        in_img_array[3][5][4] <= img[562];\
        in_img_array[3][5][5] <= img[563];\
        in_img_array[3][5][6] <= img[564];\
        in_img_array[3][5][7] <= img[565];\
        in_img_array[3][5][8] <= img[566];\
        in_img_array[3][5][9] <= img[567];\
        in_img_array[3][5][10] <= img[568];\
        in_img_array[3][5][11] <= img[569];\
        in_img_array[3][5][12] <= img[570];\
        in_img_array[3][5][13] <= img[571];\
        in_img_array[3][5][14] <= img[572];\
        in_img_array[3][5][15] <= img[573];\
        in_img_array[3][5][16] <= img[574];\
        in_img_array[3][5][17] <= img[575];\
        in_img_array[3][6][0] <= img[576];\
        in_img_array[3][6][1] <= img[577];\
        in_img_array[3][6][2] <= img[578];\
        in_img_array[3][6][3] <= img[579];\
        in_img_array[3][6][4] <= img[580];\
        in_img_array[3][6][5] <= img[581];\
        in_img_array[3][6][6] <= img[582];\
        in_img_array[3][6][7] <= img[583];\
        in_img_array[3][6][8] <= img[584];\
        in_img_array[3][6][9] <= img[585];\
        in_img_array[3][6][10] <= img[586];\
        in_img_array[3][6][11] <= img[587];\
        in_img_array[3][6][12] <= img[588];\
        in_img_array[3][6][13] <= img[589];\
        in_img_array[3][6][14] <= img[590];\
        in_img_array[3][6][15] <= img[591];\
        in_img_array[3][6][16] <= img[592];\
        in_img_array[3][6][17] <= img[593];\
        in_img_array[3][7][0] <= img[594];\
        in_img_array[3][7][1] <= img[595];\
        in_img_array[3][7][2] <= img[596];\
        in_img_array[3][7][3] <= img[597];\
        in_img_array[3][7][4] <= img[598];\
        in_img_array[3][7][5] <= img[599];\
        in_img_array[3][7][6] <= img[600];\
        in_img_array[3][7][7] <= img[601];\
        in_img_array[3][7][8] <= img[602];\
        in_img_array[3][7][9] <= img[603];\
        in_img_array[3][7][10] <= img[604];\
        in_img_array[3][7][11] <= img[605];\
        in_img_array[3][7][12] <= img[606];\
        in_img_array[3][7][13] <= img[607];\
        in_img_array[3][7][14] <= img[608];\
        in_img_array[3][7][15] <= img[609];\
        in_img_array[3][7][16] <= img[610];\
        in_img_array[3][7][17] <= img[611];\
        in_img_array[3][8][0] <= img[612];\
        in_img_array[3][8][1] <= img[613];\
        in_img_array[3][8][2] <= img[614];\
        in_img_array[3][8][3] <= img[615];\
        in_img_array[3][8][4] <= img[616];\
        in_img_array[3][8][5] <= img[617];\
        in_img_array[3][8][6] <= img[618];\
        in_img_array[3][8][7] <= img[619];\
        in_img_array[3][8][8] <= img[620];\
        in_img_array[3][8][9] <= img[621];\
        in_img_array[3][8][10] <= img[622];\
        in_img_array[3][8][11] <= img[623];\
        in_img_array[3][8][12] <= img[624];\
        in_img_array[3][8][13] <= img[625];\
        in_img_array[3][8][14] <= img[626];\
        in_img_array[3][8][15] <= img[627];\
        in_img_array[3][8][16] <= img[628];\
        in_img_array[3][8][17] <= img[629];\
        in_img_array[3][9][0] <= img[630];\
        in_img_array[3][9][1] <= img[631];\
        in_img_array[3][9][2] <= img[632];\
        in_img_array[3][9][3] <= img[633];\
        in_img_array[3][9][4] <= img[634];\
        in_img_array[3][9][5] <= img[635];\
        in_img_array[3][9][6] <= img[636];\
        in_img_array[3][9][7] <= img[637];\
        in_img_array[3][9][8] <= img[638];\
        in_img_array[3][9][9] <= img[639];\
        in_img_array[3][9][10] <= img[640];\
        in_img_array[3][9][11] <= img[641];\
        in_img_array[3][9][12] <= img[642];\
        in_img_array[3][9][13] <= img[643];\
        in_img_array[3][9][14] <= img[644];\
        in_img_array[3][9][15] <= img[645];\
        in_img_array[3][9][16] <= img[646];\
        in_img_array[3][9][17] <= img[647];\
        in_img_array[3][10][0] <= img[648];\
        in_img_array[3][10][1] <= img[649];\
        in_img_array[3][10][2] <= img[650];\
        in_img_array[3][10][3] <= img[651];\
        in_img_array[3][10][4] <= img[652];\
        in_img_array[3][10][5] <= img[653];\
        in_img_array[3][10][6] <= img[654];\
        in_img_array[3][10][7] <= img[655];\
        in_img_array[3][10][8] <= img[656];\
        in_img_array[3][10][9] <= img[657];\
        in_img_array[3][10][10] <= img[658];\
        in_img_array[3][10][11] <= img[659];\
        in_img_array[3][10][12] <= img[660];\
        in_img_array[3][10][13] <= img[661];\
        in_img_array[3][10][14] <= img[662];\
        in_img_array[3][10][15] <= img[663];\
        in_img_array[3][10][16] <= img[664];\
        in_img_array[3][10][17] <= img[665];\
        in_img_array[3][11][0] <= img[666];\
        in_img_array[3][11][1] <= img[667];\
        in_img_array[3][11][2] <= img[668];\
        in_img_array[3][11][3] <= img[669];\
        in_img_array[3][11][4] <= img[670];\
        in_img_array[3][11][5] <= img[671];\
        in_img_array[3][11][6] <= img[672];\
        in_img_array[3][11][7] <= img[673];\
        in_img_array[3][11][8] <= img[674];\
        in_img_array[3][11][9] <= img[675];\
        in_img_array[3][11][10] <= img[676];\
        in_img_array[3][11][11] <= img[677];\
        in_img_array[3][11][12] <= img[678];\
        in_img_array[3][11][13] <= img[679];\
        in_img_array[3][11][14] <= img[680];\
        in_img_array[3][11][15] <= img[681];\
        in_img_array[3][11][16] <= img[682];\
        in_img_array[3][11][17] <= img[683];\
        in_img_array[3][12][0] <= img[684];\
        in_img_array[3][12][1] <= img[685];\
        in_img_array[3][12][2] <= img[686];\
        in_img_array[3][12][3] <= img[687];\
        in_img_array[3][12][4] <= img[688];\
        in_img_array[3][12][5] <= img[689];\
        in_img_array[3][12][6] <= img[690];\
        in_img_array[3][12][7] <= img[691];\
        in_img_array[3][12][8] <= img[692];\
        in_img_array[3][12][9] <= img[693];\
        in_img_array[3][12][10] <= img[694];\
        in_img_array[3][12][11] <= img[695];\
        in_img_array[3][12][12] <= img[696];\
        in_img_array[3][12][13] <= img[697];\
        in_img_array[3][12][14] <= img[698];\
        in_img_array[3][12][15] <= img[699];\
        in_img_array[3][12][16] <= img[700];\
        in_img_array[3][12][17] <= img[701];\
        in_img_array[3][13][0] <= img[702];\
        in_img_array[3][13][1] <= img[703];\
        in_img_array[3][13][2] <= img[704];\
        in_img_array[3][13][3] <= img[705];\
        in_img_array[3][13][4] <= img[706];\
        in_img_array[3][13][5] <= img[707];\
        in_img_array[3][13][6] <= img[708];\
        in_img_array[3][13][7] <= img[709];\
        in_img_array[3][13][8] <= img[710];\
        in_img_array[3][13][9] <= img[711];\
        in_img_array[3][13][10] <= img[712];\
        in_img_array[3][13][11] <= img[713];\
        in_img_array[3][13][12] <= img[714];\
        in_img_array[3][13][13] <= img[715];\
        in_img_array[3][13][14] <= img[716];\
        in_img_array[3][13][15] <= img[717];\
        in_img_array[3][13][16] <= img[718];\
        in_img_array[3][13][17] <= img[719];\
        in_img_array[3][14][0] <= img[720];\
        in_img_array[3][14][1] <= img[721];\
        in_img_array[3][14][2] <= img[722];\
        in_img_array[3][14][3] <= img[723];\
        in_img_array[3][14][4] <= img[724];\
        in_img_array[3][14][5] <= img[725];\
        in_img_array[3][14][6] <= img[726];\
        in_img_array[3][14][7] <= img[727];\
        in_img_array[3][14][8] <= img[728];\
        in_img_array[3][14][9] <= img[729];\
        in_img_array[3][14][10] <= img[730];\
        in_img_array[3][14][11] <= img[731];\
        in_img_array[3][14][12] <= img[732];\
        in_img_array[3][14][13] <= img[733];\
        in_img_array[3][14][14] <= img[734];\
        in_img_array[3][14][15] <= img[735];\
        in_img_array[3][14][16] <= img[736];\
        in_img_array[3][14][17] <= img[737];\
        in_img_array[3][15][0] <= img[738];\
        in_img_array[3][15][1] <= img[739];\
        in_img_array[3][15][2] <= img[740];\
        in_img_array[3][15][3] <= img[741];\
        in_img_array[3][15][4] <= img[742];\
        in_img_array[3][15][5] <= img[743];\
        in_img_array[3][15][6] <= img[744];\
        in_img_array[3][15][7] <= img[745];\
        in_img_array[3][15][8] <= img[746];\
        in_img_array[3][15][9] <= img[747];\
        in_img_array[3][15][10] <= img[748];\
        in_img_array[3][15][11] <= img[749];\
        in_img_array[3][15][12] <= img[750];\
        in_img_array[3][15][13] <= img[751];\
        in_img_array[3][15][14] <= img[752];\
        in_img_array[3][15][15] <= img[753];\
        in_img_array[3][15][16] <= img[754];\
        in_img_array[3][15][17] <= img[755];\
        in_img_array[3][16][0] <= img[756];\
        in_img_array[3][16][1] <= img[757];\
        in_img_array[3][16][2] <= img[758];\
        in_img_array[3][16][3] <= img[759];\
        in_img_array[3][16][4] <= img[760];\
        in_img_array[3][16][5] <= img[761];\
        in_img_array[3][16][6] <= img[762];\
        in_img_array[3][16][7] <= img[763];\
        in_img_array[3][16][8] <= img[764];\
        in_img_array[3][16][9] <= img[765];\
        in_img_array[3][16][10] <= img[766];\
        in_img_array[3][16][11] <= img[767];\
        in_img_array[3][16][12] <= img[768];\
        in_img_array[3][16][13] <= img[769];\
        in_img_array[3][16][14] <= img[770];\
        in_img_array[3][16][15] <= img[771];\
        in_img_array[3][16][16] <= img[772];\
        in_img_array[3][16][17] <= img[773];\
        in_img_array[3][17][0] <= img[774];\
        in_img_array[3][17][1] <= img[775];\
        in_img_array[3][17][2] <= img[776];\
        in_img_array[3][17][3] <= img[777];\
        in_img_array[3][17][4] <= img[778];\
        in_img_array[3][17][5] <= img[779];\
        in_img_array[3][17][6] <= img[780];\
        in_img_array[3][17][7] <= img[781];\
        in_img_array[3][17][8] <= img[782];\
        in_img_array[3][17][9] <= img[783];\
        in_img_array[3][17][10] <= img[784];\
        in_img_array[3][17][11] <= img[785];\
        in_img_array[3][17][12] <= img[786];\
        in_img_array[3][17][13] <= img[787];\
        in_img_array[3][17][14] <= img[788];\
        in_img_array[3][17][15] <= img[789];\
        in_img_array[3][17][16] <= img[790];\
        in_img_array[3][17][17] <= img[791];\
        in_img_array[3][18][0] <= img[792];\
        in_img_array[3][18][1] <= img[793];\
        in_img_array[3][18][2] <= img[794];\
        in_img_array[3][18][3] <= img[795];\
        in_img_array[3][18][4] <= img[796];\
        in_img_array[3][18][5] <= img[797];\
        in_img_array[3][18][6] <= img[798];\
        in_img_array[3][18][7] <= img[799];\
        in_img_array[3][18][8] <= img[800];\
        in_img_array[3][18][9] <= img[801];\
        in_img_array[3][18][10] <= img[802];\
        in_img_array[3][18][11] <= img[803];\
        in_img_array[3][18][12] <= img[804];\
        in_img_array[3][18][13] <= img[805];\
        in_img_array[3][18][14] <= img[806];\
        in_img_array[3][18][15] <= img[807];\
        in_img_array[3][18][16] <= img[808];\
        in_img_array[3][18][17] <= img[809];\
        in_img_array[3][19][0] <= img[810];\
        in_img_array[3][19][1] <= img[811];\
        in_img_array[3][19][2] <= img[812];\
        in_img_array[3][19][3] <= img[813];\
        in_img_array[3][19][4] <= img[814];\
        in_img_array[3][19][5] <= img[815];\
        in_img_array[3][19][6] <= img[816];\
        in_img_array[3][19][7] <= img[817];\
        in_img_array[3][19][8] <= img[818];\
        in_img_array[3][19][9] <= img[819];\
        in_img_array[3][19][10] <= img[820];\
        in_img_array[3][19][11] <= img[821];\
        in_img_array[3][19][12] <= img[822];\
        in_img_array[3][19][13] <= img[823];\
        in_img_array[3][19][14] <= img[824];\
        in_img_array[3][19][15] <= img[825];\
        in_img_array[3][19][16] <= img[826];\
        in_img_array[3][19][17] <= img[827];\
        in_img_array[3][20][0] <= img[828];\
        in_img_array[3][20][1] <= img[829];\
        in_img_array[3][20][2] <= img[830];\
        in_img_array[3][20][3] <= img[831];\
        in_img_array[3][20][4] <= img[832];\
        in_img_array[3][20][5] <= img[833];\
        in_img_array[3][20][6] <= img[834];\
        in_img_array[3][20][7] <= img[835];\
        in_img_array[3][20][8] <= img[836];\
        in_img_array[3][20][9] <= img[837];\
        in_img_array[3][20][10] <= img[838];\
        in_img_array[3][20][11] <= img[839];\
        in_img_array[3][20][12] <= img[840];\
        in_img_array[3][20][13] <= img[841];\
        in_img_array[3][20][14] <= img[842];\
        in_img_array[3][20][15] <= img[843];\
        in_img_array[3][20][16] <= img[844];\
        in_img_array[3][20][17] <= img[845];\
        in_img_array[3][21][0] <= img[846];\
        in_img_array[3][21][1] <= img[847];\
        in_img_array[3][21][2] <= img[848];\
        in_img_array[3][21][3] <= img[849];\
        in_img_array[3][21][4] <= img[850];\
        in_img_array[3][21][5] <= img[851];\
        in_img_array[3][21][6] <= img[852];\
        in_img_array[3][21][7] <= img[853];\
        in_img_array[3][21][8] <= img[854];\
        in_img_array[3][21][9] <= img[855];\
        in_img_array[3][21][10] <= img[856];\
        in_img_array[3][21][11] <= img[857];\
        in_img_array[3][21][12] <= img[858];\
        in_img_array[3][21][13] <= img[859];\
        in_img_array[3][21][14] <= img[860];\
        in_img_array[3][21][15] <= img[861];\
        in_img_array[3][21][16] <= img[862];\
        in_img_array[3][21][17] <= img[863];\
        in_img_array[3][22][0] <= img[864];\
        in_img_array[3][22][1] <= img[865];\
        in_img_array[3][22][2] <= img[866];\
        in_img_array[3][22][3] <= img[867];\
        in_img_array[3][22][4] <= img[868];\
        in_img_array[3][22][5] <= img[869];\
        in_img_array[3][22][6] <= img[870];\
        in_img_array[3][22][7] <= img[871];\
        in_img_array[3][22][8] <= img[872];\
        in_img_array[3][22][9] <= img[873];\
        in_img_array[3][22][10] <= img[874];\
        in_img_array[3][22][11] <= img[875];\
        in_img_array[3][22][12] <= img[876];\
        in_img_array[3][22][13] <= img[877];\
        in_img_array[3][22][14] <= img[878];\
        in_img_array[3][22][15] <= img[879];\
        in_img_array[3][22][16] <= img[880];\
        in_img_array[3][22][17] <= img[881];\
        in_img_array[3][23][0] <= img[882];\
        in_img_array[3][23][1] <= img[883];\
        in_img_array[3][23][2] <= img[884];\
        in_img_array[3][23][3] <= img[885];\
        in_img_array[3][23][4] <= img[886];\
        in_img_array[3][23][5] <= img[887];\
        in_img_array[3][23][6] <= img[888];\
        in_img_array[3][23][7] <= img[889];\
        in_img_array[3][23][8] <= img[890];\
        in_img_array[3][23][9] <= img[891];\
        in_img_array[3][23][10] <= img[892];\
        in_img_array[3][23][11] <= img[893];\
        in_img_array[3][23][12] <= img[894];\
        in_img_array[3][23][13] <= img[895];\
        in_img_array[3][23][14] <= img[896];\
        in_img_array[3][23][15] <= img[897];\
        in_img_array[3][23][16] <= img[898];\
        in_img_array[3][23][17] <= img[899];\
        in_img_array[3][24][0] <= img[900];\
        in_img_array[3][24][1] <= img[901];\
        in_img_array[3][24][2] <= img[902];\
        in_img_array[3][24][3] <= img[903];\
        in_img_array[3][24][4] <= img[904];\
        in_img_array[3][24][5] <= img[905];\
        in_img_array[3][24][6] <= img[906];\
        in_img_array[3][24][7] <= img[907];\
        in_img_array[3][24][8] <= img[908];\
        in_img_array[3][24][9] <= img[909];\
        in_img_array[3][24][10] <= img[910];\
        in_img_array[3][24][11] <= img[911];\
        in_img_array[3][24][12] <= img[912];\
        in_img_array[3][24][13] <= img[913];\
        in_img_array[3][24][14] <= img[914];\
        in_img_array[3][24][15] <= img[915];\
        in_img_array[3][24][16] <= img[916];\
        in_img_array[3][24][17] <= img[917];\
        in_img_array[3][25][0] <= img[918];\
        in_img_array[3][25][1] <= img[919];\
        in_img_array[3][25][2] <= img[920];\
        in_img_array[3][25][3] <= img[921];\
        in_img_array[3][25][4] <= img[922];\
        in_img_array[3][25][5] <= img[923];\
        in_img_array[3][25][6] <= img[924];\
        in_img_array[3][25][7] <= img[925];\
        in_img_array[3][25][8] <= img[926];\
        in_img_array[3][25][9] <= img[927];\
        in_img_array[3][25][10] <= img[928];\
        in_img_array[3][25][11] <= img[929];\
        in_img_array[3][25][12] <= img[930];\
        in_img_array[3][25][13] <= img[931];\
        in_img_array[3][25][14] <= img[932];\
        in_img_array[3][25][15] <= img[933];\
        in_img_array[3][25][16] <= img[934];\
        in_img_array[3][25][17] <= img[935];\
        in_img_array[3][26][0] <= img[936];\
        in_img_array[3][26][1] <= img[937];\
        in_img_array[3][26][2] <= img[938];\
        in_img_array[3][26][3] <= img[939];\
        in_img_array[3][26][4] <= img[940];\
        in_img_array[3][26][5] <= img[941];\
        in_img_array[3][26][6] <= img[942];\
        in_img_array[3][26][7] <= img[943];\
        in_img_array[3][26][8] <= img[944];\
        in_img_array[3][26][9] <= img[945];\
        in_img_array[3][26][10] <= img[946];\
        in_img_array[3][26][11] <= img[947];\
        in_img_array[3][26][12] <= img[948];\
        in_img_array[3][26][13] <= img[949];\
        in_img_array[3][26][14] <= img[950];\
        in_img_array[3][26][15] <= img[951];\
        in_img_array[3][26][16] <= img[952];\
        in_img_array[3][26][17] <= img[953];\
        in_img_array[3][27][0] <= img[954];\
        in_img_array[3][27][1] <= img[955];\
        in_img_array[3][27][2] <= img[956];\
        in_img_array[3][27][3] <= img[957];\
        in_img_array[3][27][4] <= img[958];\
        in_img_array[3][27][5] <= img[959];\
        in_img_array[3][27][6] <= img[960];\
        in_img_array[3][27][7] <= img[961];\
        in_img_array[3][27][8] <= img[962];\
        in_img_array[3][27][9] <= img[963];\
        in_img_array[3][27][10] <= img[964];\
        in_img_array[3][27][11] <= img[965];\
        in_img_array[3][27][12] <= img[966];\
        in_img_array[3][27][13] <= img[967];\
        in_img_array[3][27][14] <= img[968];\
        in_img_array[3][27][15] <= img[969];\
        in_img_array[3][27][16] <= img[970];\
        in_img_array[3][27][17] <= img[971];\
        in_img_array[3][28][0] <= img[972];\
        in_img_array[3][28][1] <= img[973];\
        in_img_array[3][28][2] <= img[974];\
        in_img_array[3][28][3] <= img[975];\
        in_img_array[3][28][4] <= img[976];\
        in_img_array[3][28][5] <= img[977];\
        in_img_array[3][28][6] <= img[978];\
        in_img_array[3][28][7] <= img[979];\
        in_img_array[3][28][8] <= img[980];\
        in_img_array[3][28][9] <= img[981];\
        in_img_array[3][28][10] <= img[982];\
        in_img_array[3][28][11] <= img[983];\
        in_img_array[3][28][12] <= img[984];\
        in_img_array[3][28][13] <= img[985];\
        in_img_array[3][28][14] <= img[986];\
        in_img_array[3][28][15] <= img[987];\
        in_img_array[3][28][16] <= img[988];\
        in_img_array[3][28][17] <= img[989];\
        in_img_array[3][29][0] <= img[990];\
        in_img_array[3][29][1] <= img[991];\
        in_img_array[3][29][2] <= img[992];\
        in_img_array[3][29][3] <= img[993];\
        in_img_array[3][29][4] <= img[994];\
        in_img_array[3][29][5] <= img[995];\
        in_img_array[3][29][6] <= img[996];\
        in_img_array[3][29][7] <= img[997];\
        in_img_array[3][29][8] <= img[998];\
        in_img_array[3][29][9] <= img[999];\
        in_img_array[3][29][10] <= img[1000];\
        in_img_array[3][29][11] <= img[1001];\
        in_img_array[3][29][12] <= img[1002];\
        in_img_array[3][29][13] <= img[1003];\
        in_img_array[3][29][14] <= img[1004];\
        in_img_array[3][29][15] <= img[1005];\
        in_img_array[3][29][16] <= img[1006];\
        in_img_array[3][29][17] <= img[1007];\
        in_img_array[4][2][0] <= img[1008];\
        in_img_array[4][2][1] <= img[1009];\
        in_img_array[4][2][2] <= img[1010];\
        in_img_array[4][2][3] <= img[1011];\
        in_img_array[4][2][4] <= img[1012];\
        in_img_array[4][2][5] <= img[1013];\
        in_img_array[4][2][6] <= img[1014];\
        in_img_array[4][2][7] <= img[1015];\
        in_img_array[4][2][8] <= img[1016];\
        in_img_array[4][2][9] <= img[1017];\
        in_img_array[4][2][10] <= img[1018];\
        in_img_array[4][2][11] <= img[1019];\
        in_img_array[4][2][12] <= img[1020];\
        in_img_array[4][2][13] <= img[1021];\
        in_img_array[4][2][14] <= img[1022];\
        in_img_array[4][2][15] <= img[1023];\
        in_img_array[4][2][16] <= img[1024];\
        in_img_array[4][2][17] <= img[1025];\
        in_img_array[4][3][0] <= img[1026];\
        in_img_array[4][3][1] <= img[1027];\
        in_img_array[4][3][2] <= img[1028];\
        in_img_array[4][3][3] <= img[1029];\
        in_img_array[4][3][4] <= img[1030];\
        in_img_array[4][3][5] <= img[1031];\
        in_img_array[4][3][6] <= img[1032];\
        in_img_array[4][3][7] <= img[1033];\
        in_img_array[4][3][8] <= img[1034];\
        in_img_array[4][3][9] <= img[1035];\
        in_img_array[4][3][10] <= img[1036];\
        in_img_array[4][3][11] <= img[1037];\
        in_img_array[4][3][12] <= img[1038];\
        in_img_array[4][3][13] <= img[1039];\
        in_img_array[4][3][14] <= img[1040];\
        in_img_array[4][3][15] <= img[1041];\
        in_img_array[4][3][16] <= img[1042];\
        in_img_array[4][3][17] <= img[1043];\
        in_img_array[4][4][0] <= img[1044];\
        in_img_array[4][4][1] <= img[1045];\
        in_img_array[4][4][2] <= img[1046];\
        in_img_array[4][4][3] <= img[1047];\
        in_img_array[4][4][4] <= img[1048];\
        in_img_array[4][4][5] <= img[1049];\
        in_img_array[4][4][6] <= img[1050];\
        in_img_array[4][4][7] <= img[1051];\
        in_img_array[4][4][8] <= img[1052];\
        in_img_array[4][4][9] <= img[1053];\
        in_img_array[4][4][10] <= img[1054];\
        in_img_array[4][4][11] <= img[1055];\
        in_img_array[4][4][12] <= img[1056];\
        in_img_array[4][4][13] <= img[1057];\
        in_img_array[4][4][14] <= img[1058];\
        in_img_array[4][4][15] <= img[1059];\
        in_img_array[4][4][16] <= img[1060];\
        in_img_array[4][4][17] <= img[1061];\
        in_img_array[4][5][0] <= img[1062];\
        in_img_array[4][5][1] <= img[1063];\
        in_img_array[4][5][2] <= img[1064];\
        in_img_array[4][5][3] <= img[1065];\
        in_img_array[4][5][4] <= img[1066];\
        in_img_array[4][5][5] <= img[1067];\
        in_img_array[4][5][6] <= img[1068];\
        in_img_array[4][5][7] <= img[1069];\
        in_img_array[4][5][8] <= img[1070];\
        in_img_array[4][5][9] <= img[1071];\
        in_img_array[4][5][10] <= img[1072];\
        in_img_array[4][5][11] <= img[1073];\
        in_img_array[4][5][12] <= img[1074];\
        in_img_array[4][5][13] <= img[1075];\
        in_img_array[4][5][14] <= img[1076];\
        in_img_array[4][5][15] <= img[1077];\
        in_img_array[4][5][16] <= img[1078];\
        in_img_array[4][5][17] <= img[1079];\
        in_img_array[4][6][0] <= img[1080];\
        in_img_array[4][6][1] <= img[1081];\
        in_img_array[4][6][2] <= img[1082];\
        in_img_array[4][6][3] <= img[1083];\
        in_img_array[4][6][4] <= img[1084];\
        in_img_array[4][6][5] <= img[1085];\
        in_img_array[4][6][6] <= img[1086];\
        in_img_array[4][6][7] <= img[1087];\
        in_img_array[4][6][8] <= img[1088];\
        in_img_array[4][6][9] <= img[1089];\
        in_img_array[4][6][10] <= img[1090];\
        in_img_array[4][6][11] <= img[1091];\
        in_img_array[4][6][12] <= img[1092];\
        in_img_array[4][6][13] <= img[1093];\
        in_img_array[4][6][14] <= img[1094];\
        in_img_array[4][6][15] <= img[1095];\
        in_img_array[4][6][16] <= img[1096];\
        in_img_array[4][6][17] <= img[1097];\
        in_img_array[4][7][0] <= img[1098];\
        in_img_array[4][7][1] <= img[1099];\
        in_img_array[4][7][2] <= img[1100];\
        in_img_array[4][7][3] <= img[1101];\
        in_img_array[4][7][4] <= img[1102];\
        in_img_array[4][7][5] <= img[1103];\
        in_img_array[4][7][6] <= img[1104];\
        in_img_array[4][7][7] <= img[1105];\
        in_img_array[4][7][8] <= img[1106];\
        in_img_array[4][7][9] <= img[1107];\
        in_img_array[4][7][10] <= img[1108];\
        in_img_array[4][7][11] <= img[1109];\
        in_img_array[4][7][12] <= img[1110];\
        in_img_array[4][7][13] <= img[1111];\
        in_img_array[4][7][14] <= img[1112];\
        in_img_array[4][7][15] <= img[1113];\
        in_img_array[4][7][16] <= img[1114];\
        in_img_array[4][7][17] <= img[1115];\
        in_img_array[4][8][0] <= img[1116];\
        in_img_array[4][8][1] <= img[1117];\
        in_img_array[4][8][2] <= img[1118];\
        in_img_array[4][8][3] <= img[1119];\
        in_img_array[4][8][4] <= img[1120];\
        in_img_array[4][8][5] <= img[1121];\
        in_img_array[4][8][6] <= img[1122];\
        in_img_array[4][8][7] <= img[1123];\
        in_img_array[4][8][8] <= img[1124];\
        in_img_array[4][8][9] <= img[1125];\
        in_img_array[4][8][10] <= img[1126];\
        in_img_array[4][8][11] <= img[1127];\
        in_img_array[4][8][12] <= img[1128];\
        in_img_array[4][8][13] <= img[1129];\
        in_img_array[4][8][14] <= img[1130];\
        in_img_array[4][8][15] <= img[1131];\
        in_img_array[4][8][16] <= img[1132];\
        in_img_array[4][8][17] <= img[1133];\
        in_img_array[4][9][0] <= img[1134];\
        in_img_array[4][9][1] <= img[1135];\
        in_img_array[4][9][2] <= img[1136];\
        in_img_array[4][9][3] <= img[1137];\
        in_img_array[4][9][4] <= img[1138];\
        in_img_array[4][9][5] <= img[1139];\
        in_img_array[4][9][6] <= img[1140];\
        in_img_array[4][9][7] <= img[1141];\
        in_img_array[4][9][8] <= img[1142];\
        in_img_array[4][9][9] <= img[1143];\
        in_img_array[4][9][10] <= img[1144];\
        in_img_array[4][9][11] <= img[1145];\
        in_img_array[4][9][12] <= img[1146];\
        in_img_array[4][9][13] <= img[1147];\
        in_img_array[4][9][14] <= img[1148];\
        in_img_array[4][9][15] <= img[1149];\
        in_img_array[4][9][16] <= img[1150];\
        in_img_array[4][9][17] <= img[1151];\
        in_img_array[4][10][0] <= img[1152];\
        in_img_array[4][10][1] <= img[1153];\
        in_img_array[4][10][2] <= img[1154];\
        in_img_array[4][10][3] <= img[1155];\
        in_img_array[4][10][4] <= img[1156];\
        in_img_array[4][10][5] <= img[1157];\
        in_img_array[4][10][6] <= img[1158];\
        in_img_array[4][10][7] <= img[1159];\
        in_img_array[4][10][8] <= img[1160];\
        in_img_array[4][10][9] <= img[1161];\
        in_img_array[4][10][10] <= img[1162];\
        in_img_array[4][10][11] <= img[1163];\
        in_img_array[4][10][12] <= img[1164];\
        in_img_array[4][10][13] <= img[1165];\
        in_img_array[4][10][14] <= img[1166];\
        in_img_array[4][10][15] <= img[1167];\
        in_img_array[4][10][16] <= img[1168];\
        in_img_array[4][10][17] <= img[1169];\
        in_img_array[4][11][0] <= img[1170];\
        in_img_array[4][11][1] <= img[1171];\
        in_img_array[4][11][2] <= img[1172];\
        in_img_array[4][11][3] <= img[1173];\
        in_img_array[4][11][4] <= img[1174];\
        in_img_array[4][11][5] <= img[1175];\
        in_img_array[4][11][6] <= img[1176];\
        in_img_array[4][11][7] <= img[1177];\
        in_img_array[4][11][8] <= img[1178];\
        in_img_array[4][11][9] <= img[1179];\
        in_img_array[4][11][10] <= img[1180];\
        in_img_array[4][11][11] <= img[1181];\
        in_img_array[4][11][12] <= img[1182];\
        in_img_array[4][11][13] <= img[1183];\
        in_img_array[4][11][14] <= img[1184];\
        in_img_array[4][11][15] <= img[1185];\
        in_img_array[4][11][16] <= img[1186];\
        in_img_array[4][11][17] <= img[1187];\
        in_img_array[4][12][0] <= img[1188];\
        in_img_array[4][12][1] <= img[1189];\
        in_img_array[4][12][2] <= img[1190];\
        in_img_array[4][12][3] <= img[1191];\
        in_img_array[4][12][4] <= img[1192];\
        in_img_array[4][12][5] <= img[1193];\
        in_img_array[4][12][6] <= img[1194];\
        in_img_array[4][12][7] <= img[1195];\
        in_img_array[4][12][8] <= img[1196];\
        in_img_array[4][12][9] <= img[1197];\
        in_img_array[4][12][10] <= img[1198];\
        in_img_array[4][12][11] <= img[1199];\
        in_img_array[4][12][12] <= img[1200];\
        in_img_array[4][12][13] <= img[1201];\
        in_img_array[4][12][14] <= img[1202];\
        in_img_array[4][12][15] <= img[1203];\
        in_img_array[4][12][16] <= img[1204];\
        in_img_array[4][12][17] <= img[1205];\
        in_img_array[4][13][0] <= img[1206];\
        in_img_array[4][13][1] <= img[1207];\
        in_img_array[4][13][2] <= img[1208];\
        in_img_array[4][13][3] <= img[1209];\
        in_img_array[4][13][4] <= img[1210];\
        in_img_array[4][13][5] <= img[1211];\
        in_img_array[4][13][6] <= img[1212];\
        in_img_array[4][13][7] <= img[1213];\
        in_img_array[4][13][8] <= img[1214];\
        in_img_array[4][13][9] <= img[1215];\
        in_img_array[4][13][10] <= img[1216];\
        in_img_array[4][13][11] <= img[1217];\
        in_img_array[4][13][12] <= img[1218];\
        in_img_array[4][13][13] <= img[1219];\
        in_img_array[4][13][14] <= img[1220];\
        in_img_array[4][13][15] <= img[1221];\
        in_img_array[4][13][16] <= img[1222];\
        in_img_array[4][13][17] <= img[1223];\
        in_img_array[4][14][0] <= img[1224];\
        in_img_array[4][14][1] <= img[1225];\
        in_img_array[4][14][2] <= img[1226];\
        in_img_array[4][14][3] <= img[1227];\
        in_img_array[4][14][4] <= img[1228];\
        in_img_array[4][14][5] <= img[1229];\
        in_img_array[4][14][6] <= img[1230];\
        in_img_array[4][14][7] <= img[1231];\
        in_img_array[4][14][8] <= img[1232];\
        in_img_array[4][14][9] <= img[1233];\
        in_img_array[4][14][10] <= img[1234];\
        in_img_array[4][14][11] <= img[1235];\
        in_img_array[4][14][12] <= img[1236];\
        in_img_array[4][14][13] <= img[1237];\
        in_img_array[4][14][14] <= img[1238];\
        in_img_array[4][14][15] <= img[1239];\
        in_img_array[4][14][16] <= img[1240];\
        in_img_array[4][14][17] <= img[1241];\
        in_img_array[4][15][0] <= img[1242];\
        in_img_array[4][15][1] <= img[1243];\
        in_img_array[4][15][2] <= img[1244];\
        in_img_array[4][15][3] <= img[1245];\
        in_img_array[4][15][4] <= img[1246];\
        in_img_array[4][15][5] <= img[1247];\
        in_img_array[4][15][6] <= img[1248];\
        in_img_array[4][15][7] <= img[1249];\
        in_img_array[4][15][8] <= img[1250];\
        in_img_array[4][15][9] <= img[1251];\
        in_img_array[4][15][10] <= img[1252];\
        in_img_array[4][15][11] <= img[1253];\
        in_img_array[4][15][12] <= img[1254];\
        in_img_array[4][15][13] <= img[1255];\
        in_img_array[4][15][14] <= img[1256];\
        in_img_array[4][15][15] <= img[1257];\
        in_img_array[4][15][16] <= img[1258];\
        in_img_array[4][15][17] <= img[1259];\
        in_img_array[4][16][0] <= img[1260];\
        in_img_array[4][16][1] <= img[1261];\
        in_img_array[4][16][2] <= img[1262];\
        in_img_array[4][16][3] <= img[1263];\
        in_img_array[4][16][4] <= img[1264];\
        in_img_array[4][16][5] <= img[1265];\
        in_img_array[4][16][6] <= img[1266];\
        in_img_array[4][16][7] <= img[1267];\
        in_img_array[4][16][8] <= img[1268];\
        in_img_array[4][16][9] <= img[1269];\
        in_img_array[4][16][10] <= img[1270];\
        in_img_array[4][16][11] <= img[1271];\
        in_img_array[4][16][12] <= img[1272];\
        in_img_array[4][16][13] <= img[1273];\
        in_img_array[4][16][14] <= img[1274];\
        in_img_array[4][16][15] <= img[1275];\
        in_img_array[4][16][16] <= img[1276];\
        in_img_array[4][16][17] <= img[1277];\
        in_img_array[4][17][0] <= img[1278];\
        in_img_array[4][17][1] <= img[1279];\
        in_img_array[4][17][2] <= img[1280];\
        in_img_array[4][17][3] <= img[1281];\
        in_img_array[4][17][4] <= img[1282];\
        in_img_array[4][17][5] <= img[1283];\
        in_img_array[4][17][6] <= img[1284];\
        in_img_array[4][17][7] <= img[1285];\
        in_img_array[4][17][8] <= img[1286];\
        in_img_array[4][17][9] <= img[1287];\
        in_img_array[4][17][10] <= img[1288];\
        in_img_array[4][17][11] <= img[1289];\
        in_img_array[4][17][12] <= img[1290];\
        in_img_array[4][17][13] <= img[1291];\
        in_img_array[4][17][14] <= img[1292];\
        in_img_array[4][17][15] <= img[1293];\
        in_img_array[4][17][16] <= img[1294];\
        in_img_array[4][17][17] <= img[1295];\
        in_img_array[4][18][0] <= img[1296];\
        in_img_array[4][18][1] <= img[1297];\
        in_img_array[4][18][2] <= img[1298];\
        in_img_array[4][18][3] <= img[1299];\
        in_img_array[4][18][4] <= img[1300];\
        in_img_array[4][18][5] <= img[1301];\
        in_img_array[4][18][6] <= img[1302];\
        in_img_array[4][18][7] <= img[1303];\
        in_img_array[4][18][8] <= img[1304];\
        in_img_array[4][18][9] <= img[1305];\
        in_img_array[4][18][10] <= img[1306];\
        in_img_array[4][18][11] <= img[1307];\
        in_img_array[4][18][12] <= img[1308];\
        in_img_array[4][18][13] <= img[1309];\
        in_img_array[4][18][14] <= img[1310];\
        in_img_array[4][18][15] <= img[1311];\
        in_img_array[4][18][16] <= img[1312];\
        in_img_array[4][18][17] <= img[1313];\
        in_img_array[4][19][0] <= img[1314];\
        in_img_array[4][19][1] <= img[1315];\
        in_img_array[4][19][2] <= img[1316];\
        in_img_array[4][19][3] <= img[1317];\
        in_img_array[4][19][4] <= img[1318];\
        in_img_array[4][19][5] <= img[1319];\
        in_img_array[4][19][6] <= img[1320];\
        in_img_array[4][19][7] <= img[1321];\
        in_img_array[4][19][8] <= img[1322];\
        in_img_array[4][19][9] <= img[1323];\
        in_img_array[4][19][10] <= img[1324];\
        in_img_array[4][19][11] <= img[1325];\
        in_img_array[4][19][12] <= img[1326];\
        in_img_array[4][19][13] <= img[1327];\
        in_img_array[4][19][14] <= img[1328];\
        in_img_array[4][19][15] <= img[1329];\
        in_img_array[4][19][16] <= img[1330];\
        in_img_array[4][19][17] <= img[1331];\
        in_img_array[4][20][0] <= img[1332];\
        in_img_array[4][20][1] <= img[1333];\
        in_img_array[4][20][2] <= img[1334];\
        in_img_array[4][20][3] <= img[1335];\
        in_img_array[4][20][4] <= img[1336];\
        in_img_array[4][20][5] <= img[1337];\
        in_img_array[4][20][6] <= img[1338];\
        in_img_array[4][20][7] <= img[1339];\
        in_img_array[4][20][8] <= img[1340];\
        in_img_array[4][20][9] <= img[1341];\
        in_img_array[4][20][10] <= img[1342];\
        in_img_array[4][20][11] <= img[1343];\
        in_img_array[4][20][12] <= img[1344];\
        in_img_array[4][20][13] <= img[1345];\
        in_img_array[4][20][14] <= img[1346];\
        in_img_array[4][20][15] <= img[1347];\
        in_img_array[4][20][16] <= img[1348];\
        in_img_array[4][20][17] <= img[1349];\
        in_img_array[4][21][0] <= img[1350];\
        in_img_array[4][21][1] <= img[1351];\
        in_img_array[4][21][2] <= img[1352];\
        in_img_array[4][21][3] <= img[1353];\
        in_img_array[4][21][4] <= img[1354];\
        in_img_array[4][21][5] <= img[1355];\
        in_img_array[4][21][6] <= img[1356];\
        in_img_array[4][21][7] <= img[1357];\
        in_img_array[4][21][8] <= img[1358];\
        in_img_array[4][21][9] <= img[1359];\
        in_img_array[4][21][10] <= img[1360];\
        in_img_array[4][21][11] <= img[1361];\
        in_img_array[4][21][12] <= img[1362];\
        in_img_array[4][21][13] <= img[1363];\
        in_img_array[4][21][14] <= img[1364];\
        in_img_array[4][21][15] <= img[1365];\
        in_img_array[4][21][16] <= img[1366];\
        in_img_array[4][21][17] <= img[1367];\
        in_img_array[4][22][0] <= img[1368];\
        in_img_array[4][22][1] <= img[1369];\
        in_img_array[4][22][2] <= img[1370];\
        in_img_array[4][22][3] <= img[1371];\
        in_img_array[4][22][4] <= img[1372];\
        in_img_array[4][22][5] <= img[1373];\
        in_img_array[4][22][6] <= img[1374];\
        in_img_array[4][22][7] <= img[1375];\
        in_img_array[4][22][8] <= img[1376];\
        in_img_array[4][22][9] <= img[1377];\
        in_img_array[4][22][10] <= img[1378];\
        in_img_array[4][22][11] <= img[1379];\
        in_img_array[4][22][12] <= img[1380];\
        in_img_array[4][22][13] <= img[1381];\
        in_img_array[4][22][14] <= img[1382];\
        in_img_array[4][22][15] <= img[1383];\
        in_img_array[4][22][16] <= img[1384];\
        in_img_array[4][22][17] <= img[1385];\
        in_img_array[4][23][0] <= img[1386];\
        in_img_array[4][23][1] <= img[1387];\
        in_img_array[4][23][2] <= img[1388];\
        in_img_array[4][23][3] <= img[1389];\
        in_img_array[4][23][4] <= img[1390];\
        in_img_array[4][23][5] <= img[1391];\
        in_img_array[4][23][6] <= img[1392];\
        in_img_array[4][23][7] <= img[1393];\
        in_img_array[4][23][8] <= img[1394];\
        in_img_array[4][23][9] <= img[1395];\
        in_img_array[4][23][10] <= img[1396];\
        in_img_array[4][23][11] <= img[1397];\
        in_img_array[4][23][12] <= img[1398];\
        in_img_array[4][23][13] <= img[1399];\
        in_img_array[4][23][14] <= img[1400];\
        in_img_array[4][23][15] <= img[1401];\
        in_img_array[4][23][16] <= img[1402];\
        in_img_array[4][23][17] <= img[1403];\
        in_img_array[4][24][0] <= img[1404];\
        in_img_array[4][24][1] <= img[1405];\
        in_img_array[4][24][2] <= img[1406];\
        in_img_array[4][24][3] <= img[1407];\
        in_img_array[4][24][4] <= img[1408];\
        in_img_array[4][24][5] <= img[1409];\
        in_img_array[4][24][6] <= img[1410];\
        in_img_array[4][24][7] <= img[1411];\
        in_img_array[4][24][8] <= img[1412];\
        in_img_array[4][24][9] <= img[1413];\
        in_img_array[4][24][10] <= img[1414];\
        in_img_array[4][24][11] <= img[1415];\
        in_img_array[4][24][12] <= img[1416];\
        in_img_array[4][24][13] <= img[1417];\
        in_img_array[4][24][14] <= img[1418];\
        in_img_array[4][24][15] <= img[1419];\
        in_img_array[4][24][16] <= img[1420];\
        in_img_array[4][24][17] <= img[1421];\
        in_img_array[4][25][0] <= img[1422];\
        in_img_array[4][25][1] <= img[1423];\
        in_img_array[4][25][2] <= img[1424];\
        in_img_array[4][25][3] <= img[1425];\
        in_img_array[4][25][4] <= img[1426];\
        in_img_array[4][25][5] <= img[1427];\
        in_img_array[4][25][6] <= img[1428];\
        in_img_array[4][25][7] <= img[1429];\
        in_img_array[4][25][8] <= img[1430];\
        in_img_array[4][25][9] <= img[1431];\
        in_img_array[4][25][10] <= img[1432];\
        in_img_array[4][25][11] <= img[1433];\
        in_img_array[4][25][12] <= img[1434];\
        in_img_array[4][25][13] <= img[1435];\
        in_img_array[4][25][14] <= img[1436];\
        in_img_array[4][25][15] <= img[1437];\
        in_img_array[4][25][16] <= img[1438];\
        in_img_array[4][25][17] <= img[1439];\
        in_img_array[4][26][0] <= img[1440];\
        in_img_array[4][26][1] <= img[1441];\
        in_img_array[4][26][2] <= img[1442];\
        in_img_array[4][26][3] <= img[1443];\
        in_img_array[4][26][4] <= img[1444];\
        in_img_array[4][26][5] <= img[1445];\
        in_img_array[4][26][6] <= img[1446];\
        in_img_array[4][26][7] <= img[1447];\
        in_img_array[4][26][8] <= img[1448];\
        in_img_array[4][26][9] <= img[1449];\
        in_img_array[4][26][10] <= img[1450];\
        in_img_array[4][26][11] <= img[1451];\
        in_img_array[4][26][12] <= img[1452];\
        in_img_array[4][26][13] <= img[1453];\
        in_img_array[4][26][14] <= img[1454];\
        in_img_array[4][26][15] <= img[1455];\
        in_img_array[4][26][16] <= img[1456];\
        in_img_array[4][26][17] <= img[1457];\
        in_img_array[4][27][0] <= img[1458];\
        in_img_array[4][27][1] <= img[1459];\
        in_img_array[4][27][2] <= img[1460];\
        in_img_array[4][27][3] <= img[1461];\
        in_img_array[4][27][4] <= img[1462];\
        in_img_array[4][27][5] <= img[1463];\
        in_img_array[4][27][6] <= img[1464];\
        in_img_array[4][27][7] <= img[1465];\
        in_img_array[4][27][8] <= img[1466];\
        in_img_array[4][27][9] <= img[1467];\
        in_img_array[4][27][10] <= img[1468];\
        in_img_array[4][27][11] <= img[1469];\
        in_img_array[4][27][12] <= img[1470];\
        in_img_array[4][27][13] <= img[1471];\
        in_img_array[4][27][14] <= img[1472];\
        in_img_array[4][27][15] <= img[1473];\
        in_img_array[4][27][16] <= img[1474];\
        in_img_array[4][27][17] <= img[1475];\
        in_img_array[4][28][0] <= img[1476];\
        in_img_array[4][28][1] <= img[1477];\
        in_img_array[4][28][2] <= img[1478];\
        in_img_array[4][28][3] <= img[1479];\
        in_img_array[4][28][4] <= img[1480];\
        in_img_array[4][28][5] <= img[1481];\
        in_img_array[4][28][6] <= img[1482];\
        in_img_array[4][28][7] <= img[1483];\
        in_img_array[4][28][8] <= img[1484];\
        in_img_array[4][28][9] <= img[1485];\
        in_img_array[4][28][10] <= img[1486];\
        in_img_array[4][28][11] <= img[1487];\
        in_img_array[4][28][12] <= img[1488];\
        in_img_array[4][28][13] <= img[1489];\
        in_img_array[4][28][14] <= img[1490];\
        in_img_array[4][28][15] <= img[1491];\
        in_img_array[4][28][16] <= img[1492];\
        in_img_array[4][28][17] <= img[1493];\
        in_img_array[4][29][0] <= img[1494];\
        in_img_array[4][29][1] <= img[1495];\
        in_img_array[4][29][2] <= img[1496];\
        in_img_array[4][29][3] <= img[1497];\
        in_img_array[4][29][4] <= img[1498];\
        in_img_array[4][29][5] <= img[1499];\
        in_img_array[4][29][6] <= img[1500];\
        in_img_array[4][29][7] <= img[1501];\
        in_img_array[4][29][8] <= img[1502];\
        in_img_array[4][29][9] <= img[1503];\
        in_img_array[4][29][10] <= img[1504];\
        in_img_array[4][29][11] <= img[1505];\
        in_img_array[4][29][12] <= img[1506];\
        in_img_array[4][29][13] <= img[1507];\
        in_img_array[4][29][14] <= img[1508];\
        in_img_array[4][29][15] <= img[1509];\
        in_img_array[4][29][16] <= img[1510];\
        in_img_array[4][29][17] <= img[1511];\
        in_img_array[5][2][0] <= img[1512];\
        in_img_array[5][2][1] <= img[1513];\
        in_img_array[5][2][2] <= img[1514];\
        in_img_array[5][2][3] <= img[1515];\
        in_img_array[5][2][4] <= img[1516];\
        in_img_array[5][2][5] <= img[1517];\
        in_img_array[5][2][6] <= img[1518];\
        in_img_array[5][2][7] <= img[1519];\
        in_img_array[5][2][8] <= img[1520];\
        in_img_array[5][2][9] <= img[1521];\
        in_img_array[5][2][10] <= img[1522];\
        in_img_array[5][2][11] <= img[1523];\
        in_img_array[5][2][12] <= img[1524];\
        in_img_array[5][2][13] <= img[1525];\
        in_img_array[5][2][14] <= img[1526];\
        in_img_array[5][2][15] <= img[1527];\
        in_img_array[5][2][16] <= img[1528];\
        in_img_array[5][2][17] <= img[1529];\
        in_img_array[5][3][0] <= img[1530];\
        in_img_array[5][3][1] <= img[1531];\
        in_img_array[5][3][2] <= img[1532];\
        in_img_array[5][3][3] <= img[1533];\
        in_img_array[5][3][4] <= img[1534];\
        in_img_array[5][3][5] <= img[1535];\
        in_img_array[5][3][6] <= img[1536];\
        in_img_array[5][3][7] <= img[1537];\
        in_img_array[5][3][8] <= img[1538];\
        in_img_array[5][3][9] <= img[1539];\
        in_img_array[5][3][10] <= img[1540];\
        in_img_array[5][3][11] <= img[1541];\
        in_img_array[5][3][12] <= img[1542];\
        in_img_array[5][3][13] <= img[1543];\
        in_img_array[5][3][14] <= img[1544];\
        in_img_array[5][3][15] <= img[1545];\
        in_img_array[5][3][16] <= img[1546];\
        in_img_array[5][3][17] <= img[1547];\
        in_img_array[5][4][0] <= img[1548];\
        in_img_array[5][4][1] <= img[1549];\
        in_img_array[5][4][2] <= img[1550];\
        in_img_array[5][4][3] <= img[1551];\
        in_img_array[5][4][4] <= img[1552];\
        in_img_array[5][4][5] <= img[1553];\
        in_img_array[5][4][6] <= img[1554];\
        in_img_array[5][4][7] <= img[1555];\
        in_img_array[5][4][8] <= img[1556];\
        in_img_array[5][4][9] <= img[1557];\
        in_img_array[5][4][10] <= img[1558];\
        in_img_array[5][4][11] <= img[1559];\
        in_img_array[5][4][12] <= img[1560];\
        in_img_array[5][4][13] <= img[1561];\
        in_img_array[5][4][14] <= img[1562];\
        in_img_array[5][4][15] <= img[1563];\
        in_img_array[5][4][16] <= img[1564];\
        in_img_array[5][4][17] <= img[1565];\
        in_img_array[5][5][0] <= img[1566];\
        in_img_array[5][5][1] <= img[1567];\
        in_img_array[5][5][2] <= img[1568];\
        in_img_array[5][5][3] <= img[1569];\
        in_img_array[5][5][4] <= img[1570];\
        in_img_array[5][5][5] <= img[1571];\
        in_img_array[5][5][6] <= img[1572];\
        in_img_array[5][5][7] <= img[1573];\
        in_img_array[5][5][8] <= img[1574];\
        in_img_array[5][5][9] <= img[1575];\
        in_img_array[5][5][10] <= img[1576];\
        in_img_array[5][5][11] <= img[1577];\
        in_img_array[5][5][12] <= img[1578];\
        in_img_array[5][5][13] <= img[1579];\
        in_img_array[5][5][14] <= img[1580];\
        in_img_array[5][5][15] <= img[1581];\
        in_img_array[5][5][16] <= img[1582];\
        in_img_array[5][5][17] <= img[1583];\
        in_img_array[5][6][0] <= img[1584];\
        in_img_array[5][6][1] <= img[1585];\
        in_img_array[5][6][2] <= img[1586];\
        in_img_array[5][6][3] <= img[1587];\
        in_img_array[5][6][4] <= img[1588];\
        in_img_array[5][6][5] <= img[1589];\
        in_img_array[5][6][6] <= img[1590];\
        in_img_array[5][6][7] <= img[1591];\
        in_img_array[5][6][8] <= img[1592];\
        in_img_array[5][6][9] <= img[1593];\
        in_img_array[5][6][10] <= img[1594];\
        in_img_array[5][6][11] <= img[1595];\
        in_img_array[5][6][12] <= img[1596];\
        in_img_array[5][6][13] <= img[1597];\
        in_img_array[5][6][14] <= img[1598];\
        in_img_array[5][6][15] <= img[1599];\
        in_img_array[5][6][16] <= img[1600];\
        in_img_array[5][6][17] <= img[1601];\
        in_img_array[5][7][0] <= img[1602];\
        in_img_array[5][7][1] <= img[1603];\
        in_img_array[5][7][2] <= img[1604];\
        in_img_array[5][7][3] <= img[1605];\
        in_img_array[5][7][4] <= img[1606];\
        in_img_array[5][7][5] <= img[1607];\
        in_img_array[5][7][6] <= img[1608];\
        in_img_array[5][7][7] <= img[1609];\
        in_img_array[5][7][8] <= img[1610];\
        in_img_array[5][7][9] <= img[1611];\
        in_img_array[5][7][10] <= img[1612];\
        in_img_array[5][7][11] <= img[1613];\
        in_img_array[5][7][12] <= img[1614];\
        in_img_array[5][7][13] <= img[1615];\
        in_img_array[5][7][14] <= img[1616];\
        in_img_array[5][7][15] <= img[1617];\
        in_img_array[5][7][16] <= img[1618];\
        in_img_array[5][7][17] <= img[1619];\
        in_img_array[5][8][0] <= img[1620];\
        in_img_array[5][8][1] <= img[1621];\
        in_img_array[5][8][2] <= img[1622];\
        in_img_array[5][8][3] <= img[1623];\
        in_img_array[5][8][4] <= img[1624];\
        in_img_array[5][8][5] <= img[1625];\
        in_img_array[5][8][6] <= img[1626];\
        in_img_array[5][8][7] <= img[1627];\
        in_img_array[5][8][8] <= img[1628];\
        in_img_array[5][8][9] <= img[1629];\
        in_img_array[5][8][10] <= img[1630];\
        in_img_array[5][8][11] <= img[1631];\
        in_img_array[5][8][12] <= img[1632];\
        in_img_array[5][8][13] <= img[1633];\
        in_img_array[5][8][14] <= img[1634];\
        in_img_array[5][8][15] <= img[1635];\
        in_img_array[5][8][16] <= img[1636];\
        in_img_array[5][8][17] <= img[1637];\
        in_img_array[5][9][0] <= img[1638];\
        in_img_array[5][9][1] <= img[1639];\
        in_img_array[5][9][2] <= img[1640];\
        in_img_array[5][9][3] <= img[1641];\
        in_img_array[5][9][4] <= img[1642];\
        in_img_array[5][9][5] <= img[1643];\
        in_img_array[5][9][6] <= img[1644];\
        in_img_array[5][9][7] <= img[1645];\
        in_img_array[5][9][8] <= img[1646];\
        in_img_array[5][9][9] <= img[1647];\
        in_img_array[5][9][10] <= img[1648];\
        in_img_array[5][9][11] <= img[1649];\
        in_img_array[5][9][12] <= img[1650];\
        in_img_array[5][9][13] <= img[1651];\
        in_img_array[5][9][14] <= img[1652];\
        in_img_array[5][9][15] <= img[1653];\
        in_img_array[5][9][16] <= img[1654];\
        in_img_array[5][9][17] <= img[1655];\
        in_img_array[5][10][0] <= img[1656];\
        in_img_array[5][10][1] <= img[1657];\
        in_img_array[5][10][2] <= img[1658];\
        in_img_array[5][10][3] <= img[1659];\
        in_img_array[5][10][4] <= img[1660];\
        in_img_array[5][10][5] <= img[1661];\
        in_img_array[5][10][6] <= img[1662];\
        in_img_array[5][10][7] <= img[1663];\
        in_img_array[5][10][8] <= img[1664];\
        in_img_array[5][10][9] <= img[1665];\
        in_img_array[5][10][10] <= img[1666];\
        in_img_array[5][10][11] <= img[1667];\
        in_img_array[5][10][12] <= img[1668];\
        in_img_array[5][10][13] <= img[1669];\
        in_img_array[5][10][14] <= img[1670];\
        in_img_array[5][10][15] <= img[1671];\
        in_img_array[5][10][16] <= img[1672];\
        in_img_array[5][10][17] <= img[1673];\
        in_img_array[5][11][0] <= img[1674];\
        in_img_array[5][11][1] <= img[1675];\
        in_img_array[5][11][2] <= img[1676];\
        in_img_array[5][11][3] <= img[1677];\
        in_img_array[5][11][4] <= img[1678];\
        in_img_array[5][11][5] <= img[1679];\
        in_img_array[5][11][6] <= img[1680];\
        in_img_array[5][11][7] <= img[1681];\
        in_img_array[5][11][8] <= img[1682];\
        in_img_array[5][11][9] <= img[1683];\
        in_img_array[5][11][10] <= img[1684];\
        in_img_array[5][11][11] <= img[1685];\
        in_img_array[5][11][12] <= img[1686];\
        in_img_array[5][11][13] <= img[1687];\
        in_img_array[5][11][14] <= img[1688];\
        in_img_array[5][11][15] <= img[1689];\
        in_img_array[5][11][16] <= img[1690];\
        in_img_array[5][11][17] <= img[1691];\
        in_img_array[5][12][0] <= img[1692];\
        in_img_array[5][12][1] <= img[1693];\
        in_img_array[5][12][2] <= img[1694];\
        in_img_array[5][12][3] <= img[1695];\
        in_img_array[5][12][4] <= img[1696];\
        in_img_array[5][12][5] <= img[1697];\
        in_img_array[5][12][6] <= img[1698];\
        in_img_array[5][12][7] <= img[1699];\
        in_img_array[5][12][8] <= img[1700];\
        in_img_array[5][12][9] <= img[1701];\
        in_img_array[5][12][10] <= img[1702];\
        in_img_array[5][12][11] <= img[1703];\
        in_img_array[5][12][12] <= img[1704];\
        in_img_array[5][12][13] <= img[1705];\
        in_img_array[5][12][14] <= img[1706];\
        in_img_array[5][12][15] <= img[1707];\
        in_img_array[5][12][16] <= img[1708];\
        in_img_array[5][12][17] <= img[1709];\
        in_img_array[5][13][0] <= img[1710];\
        in_img_array[5][13][1] <= img[1711];\
        in_img_array[5][13][2] <= img[1712];\
        in_img_array[5][13][3] <= img[1713];\
        in_img_array[5][13][4] <= img[1714];\
        in_img_array[5][13][5] <= img[1715];\
        in_img_array[5][13][6] <= img[1716];\
        in_img_array[5][13][7] <= img[1717];\
        in_img_array[5][13][8] <= img[1718];\
        in_img_array[5][13][9] <= img[1719];\
        in_img_array[5][13][10] <= img[1720];\
        in_img_array[5][13][11] <= img[1721];\
        in_img_array[5][13][12] <= img[1722];\
        in_img_array[5][13][13] <= img[1723];\
        in_img_array[5][13][14] <= img[1724];\
        in_img_array[5][13][15] <= img[1725];\
        in_img_array[5][13][16] <= img[1726];\
        in_img_array[5][13][17] <= img[1727];\
        in_img_array[5][14][0] <= img[1728];\
        in_img_array[5][14][1] <= img[1729];\
        in_img_array[5][14][2] <= img[1730];\
        in_img_array[5][14][3] <= img[1731];\
        in_img_array[5][14][4] <= img[1732];\
        in_img_array[5][14][5] <= img[1733];\
        in_img_array[5][14][6] <= img[1734];\
        in_img_array[5][14][7] <= img[1735];\
        in_img_array[5][14][8] <= img[1736];\
        in_img_array[5][14][9] <= img[1737];\
        in_img_array[5][14][10] <= img[1738];\
        in_img_array[5][14][11] <= img[1739];\
        in_img_array[5][14][12] <= img[1740];\
        in_img_array[5][14][13] <= img[1741];\
        in_img_array[5][14][14] <= img[1742];\
        in_img_array[5][14][15] <= img[1743];\
        in_img_array[5][14][16] <= img[1744];\
        in_img_array[5][14][17] <= img[1745];\
        in_img_array[5][15][0] <= img[1746];\
        in_img_array[5][15][1] <= img[1747];\
        in_img_array[5][15][2] <= img[1748];\
        in_img_array[5][15][3] <= img[1749];\
        in_img_array[5][15][4] <= img[1750];\
        in_img_array[5][15][5] <= img[1751];\
        in_img_array[5][15][6] <= img[1752];\
        in_img_array[5][15][7] <= img[1753];\
        in_img_array[5][15][8] <= img[1754];\
        in_img_array[5][15][9] <= img[1755];\
        in_img_array[5][15][10] <= img[1756];\
        in_img_array[5][15][11] <= img[1757];\
        in_img_array[5][15][12] <= img[1758];\
        in_img_array[5][15][13] <= img[1759];\
        in_img_array[5][15][14] <= img[1760];\
        in_img_array[5][15][15] <= img[1761];\
        in_img_array[5][15][16] <= img[1762];\
        in_img_array[5][15][17] <= img[1763];\
        in_img_array[5][16][0] <= img[1764];\
        in_img_array[5][16][1] <= img[1765];\
        in_img_array[5][16][2] <= img[1766];\
        in_img_array[5][16][3] <= img[1767];\
        in_img_array[5][16][4] <= img[1768];\
        in_img_array[5][16][5] <= img[1769];\
        in_img_array[5][16][6] <= img[1770];\
        in_img_array[5][16][7] <= img[1771];\
        in_img_array[5][16][8] <= img[1772];\
        in_img_array[5][16][9] <= img[1773];\
        in_img_array[5][16][10] <= img[1774];\
        in_img_array[5][16][11] <= img[1775];\
        in_img_array[5][16][12] <= img[1776];\
        in_img_array[5][16][13] <= img[1777];\
        in_img_array[5][16][14] <= img[1778];\
        in_img_array[5][16][15] <= img[1779];\
        in_img_array[5][16][16] <= img[1780];\
        in_img_array[5][16][17] <= img[1781];\
        in_img_array[5][17][0] <= img[1782];\
        in_img_array[5][17][1] <= img[1783];\
        in_img_array[5][17][2] <= img[1784];\
        in_img_array[5][17][3] <= img[1785];\
        in_img_array[5][17][4] <= img[1786];\
        in_img_array[5][17][5] <= img[1787];\
        in_img_array[5][17][6] <= img[1788];\
        in_img_array[5][17][7] <= img[1789];\
        in_img_array[5][17][8] <= img[1790];\
        in_img_array[5][17][9] <= img[1791];\
        in_img_array[5][17][10] <= img[1792];\
        in_img_array[5][17][11] <= img[1793];\
        in_img_array[5][17][12] <= img[1794];\
        in_img_array[5][17][13] <= img[1795];\
        in_img_array[5][17][14] <= img[1796];\
        in_img_array[5][17][15] <= img[1797];\
        in_img_array[5][17][16] <= img[1798];\
        in_img_array[5][17][17] <= img[1799];\
        in_img_array[5][18][0] <= img[1800];\
        in_img_array[5][18][1] <= img[1801];\
        in_img_array[5][18][2] <= img[1802];\
        in_img_array[5][18][3] <= img[1803];\
        in_img_array[5][18][4] <= img[1804];\
        in_img_array[5][18][5] <= img[1805];\
        in_img_array[5][18][6] <= img[1806];\
        in_img_array[5][18][7] <= img[1807];\
        in_img_array[5][18][8] <= img[1808];\
        in_img_array[5][18][9] <= img[1809];\
        in_img_array[5][18][10] <= img[1810];\
        in_img_array[5][18][11] <= img[1811];\
        in_img_array[5][18][12] <= img[1812];\
        in_img_array[5][18][13] <= img[1813];\
        in_img_array[5][18][14] <= img[1814];\
        in_img_array[5][18][15] <= img[1815];\
        in_img_array[5][18][16] <= img[1816];\
        in_img_array[5][18][17] <= img[1817];\
        in_img_array[5][19][0] <= img[1818];\
        in_img_array[5][19][1] <= img[1819];\
        in_img_array[5][19][2] <= img[1820];\
        in_img_array[5][19][3] <= img[1821];\
        in_img_array[5][19][4] <= img[1822];\
        in_img_array[5][19][5] <= img[1823];\
        in_img_array[5][19][6] <= img[1824];\
        in_img_array[5][19][7] <= img[1825];\
        in_img_array[5][19][8] <= img[1826];\
        in_img_array[5][19][9] <= img[1827];\
        in_img_array[5][19][10] <= img[1828];\
        in_img_array[5][19][11] <= img[1829];\
        in_img_array[5][19][12] <= img[1830];\
        in_img_array[5][19][13] <= img[1831];\
        in_img_array[5][19][14] <= img[1832];\
        in_img_array[5][19][15] <= img[1833];\
        in_img_array[5][19][16] <= img[1834];\
        in_img_array[5][19][17] <= img[1835];\
        in_img_array[5][20][0] <= img[1836];\
        in_img_array[5][20][1] <= img[1837];\
        in_img_array[5][20][2] <= img[1838];\
        in_img_array[5][20][3] <= img[1839];\
        in_img_array[5][20][4] <= img[1840];\
        in_img_array[5][20][5] <= img[1841];\
        in_img_array[5][20][6] <= img[1842];\
        in_img_array[5][20][7] <= img[1843];\
        in_img_array[5][20][8] <= img[1844];\
        in_img_array[5][20][9] <= img[1845];\
        in_img_array[5][20][10] <= img[1846];\
        in_img_array[5][20][11] <= img[1847];\
        in_img_array[5][20][12] <= img[1848];\
        in_img_array[5][20][13] <= img[1849];\
        in_img_array[5][20][14] <= img[1850];\
        in_img_array[5][20][15] <= img[1851];\
        in_img_array[5][20][16] <= img[1852];\
        in_img_array[5][20][17] <= img[1853];\
        in_img_array[5][21][0] <= img[1854];\
        in_img_array[5][21][1] <= img[1855];\
        in_img_array[5][21][2] <= img[1856];\
        in_img_array[5][21][3] <= img[1857];\
        in_img_array[5][21][4] <= img[1858];\
        in_img_array[5][21][5] <= img[1859];\
        in_img_array[5][21][6] <= img[1860];\
        in_img_array[5][21][7] <= img[1861];\
        in_img_array[5][21][8] <= img[1862];\
        in_img_array[5][21][9] <= img[1863];\
        in_img_array[5][21][10] <= img[1864];\
        in_img_array[5][21][11] <= img[1865];\
        in_img_array[5][21][12] <= img[1866];\
        in_img_array[5][21][13] <= img[1867];\
        in_img_array[5][21][14] <= img[1868];\
        in_img_array[5][21][15] <= img[1869];\
        in_img_array[5][21][16] <= img[1870];\
        in_img_array[5][21][17] <= img[1871];\
        in_img_array[5][22][0] <= img[1872];\
        in_img_array[5][22][1] <= img[1873];\
        in_img_array[5][22][2] <= img[1874];\
        in_img_array[5][22][3] <= img[1875];\
        in_img_array[5][22][4] <= img[1876];\
        in_img_array[5][22][5] <= img[1877];\
        in_img_array[5][22][6] <= img[1878];\
        in_img_array[5][22][7] <= img[1879];\
        in_img_array[5][22][8] <= img[1880];\
        in_img_array[5][22][9] <= img[1881];\
        in_img_array[5][22][10] <= img[1882];\
        in_img_array[5][22][11] <= img[1883];\
        in_img_array[5][22][12] <= img[1884];\
        in_img_array[5][22][13] <= img[1885];\
        in_img_array[5][22][14] <= img[1886];\
        in_img_array[5][22][15] <= img[1887];\
        in_img_array[5][22][16] <= img[1888];\
        in_img_array[5][22][17] <= img[1889];\
        in_img_array[5][23][0] <= img[1890];\
        in_img_array[5][23][1] <= img[1891];\
        in_img_array[5][23][2] <= img[1892];\
        in_img_array[5][23][3] <= img[1893];\
        in_img_array[5][23][4] <= img[1894];\
        in_img_array[5][23][5] <= img[1895];\
        in_img_array[5][23][6] <= img[1896];\
        in_img_array[5][23][7] <= img[1897];\
        in_img_array[5][23][8] <= img[1898];\
        in_img_array[5][23][9] <= img[1899];\
        in_img_array[5][23][10] <= img[1900];\
        in_img_array[5][23][11] <= img[1901];\
        in_img_array[5][23][12] <= img[1902];\
        in_img_array[5][23][13] <= img[1903];\
        in_img_array[5][23][14] <= img[1904];\
        in_img_array[5][23][15] <= img[1905];\
        in_img_array[5][23][16] <= img[1906];\
        in_img_array[5][23][17] <= img[1907];\
        in_img_array[5][24][0] <= img[1908];\
        in_img_array[5][24][1] <= img[1909];\
        in_img_array[5][24][2] <= img[1910];\
        in_img_array[5][24][3] <= img[1911];\
        in_img_array[5][24][4] <= img[1912];\
        in_img_array[5][24][5] <= img[1913];\
        in_img_array[5][24][6] <= img[1914];\
        in_img_array[5][24][7] <= img[1915];\
        in_img_array[5][24][8] <= img[1916];\
        in_img_array[5][24][9] <= img[1917];\
        in_img_array[5][24][10] <= img[1918];\
        in_img_array[5][24][11] <= img[1919];\
        in_img_array[5][24][12] <= img[1920];\
        in_img_array[5][24][13] <= img[1921];\
        in_img_array[5][24][14] <= img[1922];\
        in_img_array[5][24][15] <= img[1923];\
        in_img_array[5][24][16] <= img[1924];\
        in_img_array[5][24][17] <= img[1925];\
        in_img_array[5][25][0] <= img[1926];\
        in_img_array[5][25][1] <= img[1927];\
        in_img_array[5][25][2] <= img[1928];\
        in_img_array[5][25][3] <= img[1929];\
        in_img_array[5][25][4] <= img[1930];\
        in_img_array[5][25][5] <= img[1931];\
        in_img_array[5][25][6] <= img[1932];\
        in_img_array[5][25][7] <= img[1933];\
        in_img_array[5][25][8] <= img[1934];\
        in_img_array[5][25][9] <= img[1935];\
        in_img_array[5][25][10] <= img[1936];\
        in_img_array[5][25][11] <= img[1937];\
        in_img_array[5][25][12] <= img[1938];\
        in_img_array[5][25][13] <= img[1939];\
        in_img_array[5][25][14] <= img[1940];\
        in_img_array[5][25][15] <= img[1941];\
        in_img_array[5][25][16] <= img[1942];\
        in_img_array[5][25][17] <= img[1943];\
        in_img_array[5][26][0] <= img[1944];\
        in_img_array[5][26][1] <= img[1945];\
        in_img_array[5][26][2] <= img[1946];\
        in_img_array[5][26][3] <= img[1947];\
        in_img_array[5][26][4] <= img[1948];\
        in_img_array[5][26][5] <= img[1949];\
        in_img_array[5][26][6] <= img[1950];\
        in_img_array[5][26][7] <= img[1951];\
        in_img_array[5][26][8] <= img[1952];\
        in_img_array[5][26][9] <= img[1953];\
        in_img_array[5][26][10] <= img[1954];\
        in_img_array[5][26][11] <= img[1955];\
        in_img_array[5][26][12] <= img[1956];\
        in_img_array[5][26][13] <= img[1957];\
        in_img_array[5][26][14] <= img[1958];\
        in_img_array[5][26][15] <= img[1959];\
        in_img_array[5][26][16] <= img[1960];\
        in_img_array[5][26][17] <= img[1961];\
        in_img_array[5][27][0] <= img[1962];\
        in_img_array[5][27][1] <= img[1963];\
        in_img_array[5][27][2] <= img[1964];\
        in_img_array[5][27][3] <= img[1965];\
        in_img_array[5][27][4] <= img[1966];\
        in_img_array[5][27][5] <= img[1967];\
        in_img_array[5][27][6] <= img[1968];\
        in_img_array[5][27][7] <= img[1969];\
        in_img_array[5][27][8] <= img[1970];\
        in_img_array[5][27][9] <= img[1971];\
        in_img_array[5][27][10] <= img[1972];\
        in_img_array[5][27][11] <= img[1973];\
        in_img_array[5][27][12] <= img[1974];\
        in_img_array[5][27][13] <= img[1975];\
        in_img_array[5][27][14] <= img[1976];\
        in_img_array[5][27][15] <= img[1977];\
        in_img_array[5][27][16] <= img[1978];\
        in_img_array[5][27][17] <= img[1979];\
        in_img_array[5][28][0] <= img[1980];\
        in_img_array[5][28][1] <= img[1981];\
        in_img_array[5][28][2] <= img[1982];\
        in_img_array[5][28][3] <= img[1983];\
        in_img_array[5][28][4] <= img[1984];\
        in_img_array[5][28][5] <= img[1985];\
        in_img_array[5][28][6] <= img[1986];\
        in_img_array[5][28][7] <= img[1987];\
        in_img_array[5][28][8] <= img[1988];\
        in_img_array[5][28][9] <= img[1989];\
        in_img_array[5][28][10] <= img[1990];\
        in_img_array[5][28][11] <= img[1991];\
        in_img_array[5][28][12] <= img[1992];\
        in_img_array[5][28][13] <= img[1993];\
        in_img_array[5][28][14] <= img[1994];\
        in_img_array[5][28][15] <= img[1995];\
        in_img_array[5][28][16] <= img[1996];\
        in_img_array[5][28][17] <= img[1997];\
        in_img_array[5][29][0] <= img[1998];\
        in_img_array[5][29][1] <= img[1999];\
        in_img_array[5][29][2] <= img[2000];\
        in_img_array[5][29][3] <= img[2001];\
        in_img_array[5][29][4] <= img[2002];\
        in_img_array[5][29][5] <= img[2003];\
        in_img_array[5][29][6] <= img[2004];\
        in_img_array[5][29][7] <= img[2005];\
        in_img_array[5][29][8] <= img[2006];\
        in_img_array[5][29][9] <= img[2007];\
        in_img_array[5][29][10] <= img[2008];\
        in_img_array[5][29][11] <= img[2009];\
        in_img_array[5][29][12] <= img[2010];\
        in_img_array[5][29][13] <= img[2011];\
        in_img_array[5][29][14] <= img[2012];\
        in_img_array[5][29][15] <= img[2013];\
        in_img_array[5][29][16] <= img[2014];\
        in_img_array[5][29][17] <= img[2015];\
        in_img_array[6][2][0] <= img[2016];\
        in_img_array[6][2][1] <= img[2017];\
        in_img_array[6][2][2] <= img[2018];\
        in_img_array[6][2][3] <= img[2019];\
        in_img_array[6][2][4] <= img[2020];\
        in_img_array[6][2][5] <= img[2021];\
        in_img_array[6][2][6] <= img[2022];\
        in_img_array[6][2][7] <= img[2023];\
        in_img_array[6][2][8] <= img[2024];\
        in_img_array[6][2][9] <= img[2025];\
        in_img_array[6][2][10] <= img[2026];\
        in_img_array[6][2][11] <= img[2027];\
        in_img_array[6][2][12] <= img[2028];\
        in_img_array[6][2][13] <= img[2029];\
        in_img_array[6][2][14] <= img[2030];\
        in_img_array[6][2][15] <= img[2031];\
        in_img_array[6][2][16] <= img[2032];\
        in_img_array[6][2][17] <= img[2033];\
        in_img_array[6][3][0] <= img[2034];\
        in_img_array[6][3][1] <= img[2035];\
        in_img_array[6][3][2] <= img[2036];\
        in_img_array[6][3][3] <= img[2037];\
        in_img_array[6][3][4] <= img[2038];\
        in_img_array[6][3][5] <= img[2039];\
        in_img_array[6][3][6] <= img[2040];\
        in_img_array[6][3][7] <= img[2041];\
        in_img_array[6][3][8] <= img[2042];\
        in_img_array[6][3][9] <= img[2043];\
        in_img_array[6][3][10] <= img[2044];\
        in_img_array[6][3][11] <= img[2045];\
        in_img_array[6][3][12] <= img[2046];\
        in_img_array[6][3][13] <= img[2047];\
        in_img_array[6][3][14] <= img[2048];\
        in_img_array[6][3][15] <= img[2049];\
        in_img_array[6][3][16] <= img[2050];\
        in_img_array[6][3][17] <= img[2051];\
        in_img_array[6][4][0] <= img[2052];\
        in_img_array[6][4][1] <= img[2053];\
        in_img_array[6][4][2] <= img[2054];\
        in_img_array[6][4][3] <= img[2055];\
        in_img_array[6][4][4] <= img[2056];\
        in_img_array[6][4][5] <= img[2057];\
        in_img_array[6][4][6] <= img[2058];\
        in_img_array[6][4][7] <= img[2059];\
        in_img_array[6][4][8] <= img[2060];\
        in_img_array[6][4][9] <= img[2061];\
        in_img_array[6][4][10] <= img[2062];\
        in_img_array[6][4][11] <= img[2063];\
        in_img_array[6][4][12] <= img[2064];\
        in_img_array[6][4][13] <= img[2065];\
        in_img_array[6][4][14] <= img[2066];\
        in_img_array[6][4][15] <= img[2067];\
        in_img_array[6][4][16] <= img[2068];\
        in_img_array[6][4][17] <= img[2069];\
        in_img_array[6][5][0] <= img[2070];\
        in_img_array[6][5][1] <= img[2071];\
        in_img_array[6][5][2] <= img[2072];\
        in_img_array[6][5][3] <= img[2073];\
        in_img_array[6][5][4] <= img[2074];\
        in_img_array[6][5][5] <= img[2075];\
        in_img_array[6][5][6] <= img[2076];\
        in_img_array[6][5][7] <= img[2077];\
        in_img_array[6][5][8] <= img[2078];\
        in_img_array[6][5][9] <= img[2079];\
        in_img_array[6][5][10] <= img[2080];\
        in_img_array[6][5][11] <= img[2081];\
        in_img_array[6][5][12] <= img[2082];\
        in_img_array[6][5][13] <= img[2083];\
        in_img_array[6][5][14] <= img[2084];\
        in_img_array[6][5][15] <= img[2085];\
        in_img_array[6][5][16] <= img[2086];\
        in_img_array[6][5][17] <= img[2087];\
        in_img_array[6][6][0] <= img[2088];\
        in_img_array[6][6][1] <= img[2089];\
        in_img_array[6][6][2] <= img[2090];\
        in_img_array[6][6][3] <= img[2091];\
        in_img_array[6][6][4] <= img[2092];\
        in_img_array[6][6][5] <= img[2093];\
        in_img_array[6][6][6] <= img[2094];\
        in_img_array[6][6][7] <= img[2095];\
        in_img_array[6][6][8] <= img[2096];\
        in_img_array[6][6][9] <= img[2097];\
        in_img_array[6][6][10] <= img[2098];\
        in_img_array[6][6][11] <= img[2099];\
        in_img_array[6][6][12] <= img[2100];\
        in_img_array[6][6][13] <= img[2101];\
        in_img_array[6][6][14] <= img[2102];\
        in_img_array[6][6][15] <= img[2103];\
        in_img_array[6][6][16] <= img[2104];\
        in_img_array[6][6][17] <= img[2105];\
        in_img_array[6][7][0] <= img[2106];\
        in_img_array[6][7][1] <= img[2107];\
        in_img_array[6][7][2] <= img[2108];\
        in_img_array[6][7][3] <= img[2109];\
        in_img_array[6][7][4] <= img[2110];\
        in_img_array[6][7][5] <= img[2111];\
        in_img_array[6][7][6] <= img[2112];\
        in_img_array[6][7][7] <= img[2113];\
        in_img_array[6][7][8] <= img[2114];\
        in_img_array[6][7][9] <= img[2115];\
        in_img_array[6][7][10] <= img[2116];\
        in_img_array[6][7][11] <= img[2117];\
        in_img_array[6][7][12] <= img[2118];\
        in_img_array[6][7][13] <= img[2119];\
        in_img_array[6][7][14] <= img[2120];\
        in_img_array[6][7][15] <= img[2121];\
        in_img_array[6][7][16] <= img[2122];\
        in_img_array[6][7][17] <= img[2123];\
        in_img_array[6][8][0] <= img[2124];\
        in_img_array[6][8][1] <= img[2125];\
        in_img_array[6][8][2] <= img[2126];\
        in_img_array[6][8][3] <= img[2127];\
        in_img_array[6][8][4] <= img[2128];\
        in_img_array[6][8][5] <= img[2129];\
        in_img_array[6][8][6] <= img[2130];\
        in_img_array[6][8][7] <= img[2131];\
        in_img_array[6][8][8] <= img[2132];\
        in_img_array[6][8][9] <= img[2133];\
        in_img_array[6][8][10] <= img[2134];\
        in_img_array[6][8][11] <= img[2135];\
        in_img_array[6][8][12] <= img[2136];\
        in_img_array[6][8][13] <= img[2137];\
        in_img_array[6][8][14] <= img[2138];\
        in_img_array[6][8][15] <= img[2139];\
        in_img_array[6][8][16] <= img[2140];\
        in_img_array[6][8][17] <= img[2141];\
        in_img_array[6][9][0] <= img[2142];\
        in_img_array[6][9][1] <= img[2143];\
        in_img_array[6][9][2] <= img[2144];\
        in_img_array[6][9][3] <= img[2145];\
        in_img_array[6][9][4] <= img[2146];\
        in_img_array[6][9][5] <= img[2147];\
        in_img_array[6][9][6] <= img[2148];\
        in_img_array[6][9][7] <= img[2149];\
        in_img_array[6][9][8] <= img[2150];\
        in_img_array[6][9][9] <= img[2151];\
        in_img_array[6][9][10] <= img[2152];\
        in_img_array[6][9][11] <= img[2153];\
        in_img_array[6][9][12] <= img[2154];\
        in_img_array[6][9][13] <= img[2155];\
        in_img_array[6][9][14] <= img[2156];\
        in_img_array[6][9][15] <= img[2157];\
        in_img_array[6][9][16] <= img[2158];\
        in_img_array[6][9][17] <= img[2159];\
        in_img_array[6][10][0] <= img[2160];\
        in_img_array[6][10][1] <= img[2161];\
        in_img_array[6][10][2] <= img[2162];\
        in_img_array[6][10][3] <= img[2163];\
        in_img_array[6][10][4] <= img[2164];\
        in_img_array[6][10][5] <= img[2165];\
        in_img_array[6][10][6] <= img[2166];\
        in_img_array[6][10][7] <= img[2167];\
        in_img_array[6][10][8] <= img[2168];\
        in_img_array[6][10][9] <= img[2169];\
        in_img_array[6][10][10] <= img[2170];\
        in_img_array[6][10][11] <= img[2171];\
        in_img_array[6][10][12] <= img[2172];\
        in_img_array[6][10][13] <= img[2173];\
        in_img_array[6][10][14] <= img[2174];\
        in_img_array[6][10][15] <= img[2175];\
        in_img_array[6][10][16] <= img[2176];\
        in_img_array[6][10][17] <= img[2177];\
        in_img_array[6][11][0] <= img[2178];\
        in_img_array[6][11][1] <= img[2179];\
        in_img_array[6][11][2] <= img[2180];\
        in_img_array[6][11][3] <= img[2181];\
        in_img_array[6][11][4] <= img[2182];\
        in_img_array[6][11][5] <= img[2183];\
        in_img_array[6][11][6] <= img[2184];\
        in_img_array[6][11][7] <= img[2185];\
        in_img_array[6][11][8] <= img[2186];\
        in_img_array[6][11][9] <= img[2187];\
        in_img_array[6][11][10] <= img[2188];\
        in_img_array[6][11][11] <= img[2189];\
        in_img_array[6][11][12] <= img[2190];\
        in_img_array[6][11][13] <= img[2191];\
        in_img_array[6][11][14] <= img[2192];\
        in_img_array[6][11][15] <= img[2193];\
        in_img_array[6][11][16] <= img[2194];\
        in_img_array[6][11][17] <= img[2195];\
        in_img_array[6][12][0] <= img[2196];\
        in_img_array[6][12][1] <= img[2197];\
        in_img_array[6][12][2] <= img[2198];\
        in_img_array[6][12][3] <= img[2199];\
        in_img_array[6][12][4] <= img[2200];\
        in_img_array[6][12][5] <= img[2201];\
        in_img_array[6][12][6] <= img[2202];\
        in_img_array[6][12][7] <= img[2203];\
        in_img_array[6][12][8] <= img[2204];\
        in_img_array[6][12][9] <= img[2205];\
        in_img_array[6][12][10] <= img[2206];\
        in_img_array[6][12][11] <= img[2207];\
        in_img_array[6][12][12] <= img[2208];\
        in_img_array[6][12][13] <= img[2209];\
        in_img_array[6][12][14] <= img[2210];\
        in_img_array[6][12][15] <= img[2211];\
        in_img_array[6][12][16] <= img[2212];\
        in_img_array[6][12][17] <= img[2213];\
        in_img_array[6][13][0] <= img[2214];\
        in_img_array[6][13][1] <= img[2215];\
        in_img_array[6][13][2] <= img[2216];\
        in_img_array[6][13][3] <= img[2217];\
        in_img_array[6][13][4] <= img[2218];\
        in_img_array[6][13][5] <= img[2219];\
        in_img_array[6][13][6] <= img[2220];\
        in_img_array[6][13][7] <= img[2221];\
        in_img_array[6][13][8] <= img[2222];\
        in_img_array[6][13][9] <= img[2223];\
        in_img_array[6][13][10] <= img[2224];\
        in_img_array[6][13][11] <= img[2225];\
        in_img_array[6][13][12] <= img[2226];\
        in_img_array[6][13][13] <= img[2227];\
        in_img_array[6][13][14] <= img[2228];\
        in_img_array[6][13][15] <= img[2229];\
        in_img_array[6][13][16] <= img[2230];\
        in_img_array[6][13][17] <= img[2231];\
        in_img_array[6][14][0] <= img[2232];\
        in_img_array[6][14][1] <= img[2233];\
        in_img_array[6][14][2] <= img[2234];\
        in_img_array[6][14][3] <= img[2235];\
        in_img_array[6][14][4] <= img[2236];\
        in_img_array[6][14][5] <= img[2237];\
        in_img_array[6][14][6] <= img[2238];\
        in_img_array[6][14][7] <= img[2239];\
        in_img_array[6][14][8] <= img[2240];\
        in_img_array[6][14][9] <= img[2241];\
        in_img_array[6][14][10] <= img[2242];\
        in_img_array[6][14][11] <= img[2243];\
        in_img_array[6][14][12] <= img[2244];\
        in_img_array[6][14][13] <= img[2245];\
        in_img_array[6][14][14] <= img[2246];\
        in_img_array[6][14][15] <= img[2247];\
        in_img_array[6][14][16] <= img[2248];\
        in_img_array[6][14][17] <= img[2249];\
        in_img_array[6][15][0] <= img[2250];\
        in_img_array[6][15][1] <= img[2251];\
        in_img_array[6][15][2] <= img[2252];\
        in_img_array[6][15][3] <= img[2253];\
        in_img_array[6][15][4] <= img[2254];\
        in_img_array[6][15][5] <= img[2255];\
        in_img_array[6][15][6] <= img[2256];\
        in_img_array[6][15][7] <= img[2257];\
        in_img_array[6][15][8] <= img[2258];\
        in_img_array[6][15][9] <= img[2259];\
        in_img_array[6][15][10] <= img[2260];\
        in_img_array[6][15][11] <= img[2261];\
        in_img_array[6][15][12] <= img[2262];\
        in_img_array[6][15][13] <= img[2263];\
        in_img_array[6][15][14] <= img[2264];\
        in_img_array[6][15][15] <= img[2265];\
        in_img_array[6][15][16] <= img[2266];\
        in_img_array[6][15][17] <= img[2267];\
        in_img_array[6][16][0] <= img[2268];\
        in_img_array[6][16][1] <= img[2269];\
        in_img_array[6][16][2] <= img[2270];\
        in_img_array[6][16][3] <= img[2271];\
        in_img_array[6][16][4] <= img[2272];\
        in_img_array[6][16][5] <= img[2273];\
        in_img_array[6][16][6] <= img[2274];\
        in_img_array[6][16][7] <= img[2275];\
        in_img_array[6][16][8] <= img[2276];\
        in_img_array[6][16][9] <= img[2277];\
        in_img_array[6][16][10] <= img[2278];\
        in_img_array[6][16][11] <= img[2279];\
        in_img_array[6][16][12] <= img[2280];\
        in_img_array[6][16][13] <= img[2281];\
        in_img_array[6][16][14] <= img[2282];\
        in_img_array[6][16][15] <= img[2283];\
        in_img_array[6][16][16] <= img[2284];\
        in_img_array[6][16][17] <= img[2285];\
        in_img_array[6][17][0] <= img[2286];\
        in_img_array[6][17][1] <= img[2287];\
        in_img_array[6][17][2] <= img[2288];\
        in_img_array[6][17][3] <= img[2289];\
        in_img_array[6][17][4] <= img[2290];\
        in_img_array[6][17][5] <= img[2291];\
        in_img_array[6][17][6] <= img[2292];\
        in_img_array[6][17][7] <= img[2293];\
        in_img_array[6][17][8] <= img[2294];\
        in_img_array[6][17][9] <= img[2295];\
        in_img_array[6][17][10] <= img[2296];\
        in_img_array[6][17][11] <= img[2297];\
        in_img_array[6][17][12] <= img[2298];\
        in_img_array[6][17][13] <= img[2299];\
        in_img_array[6][17][14] <= img[2300];\
        in_img_array[6][17][15] <= img[2301];\
        in_img_array[6][17][16] <= img[2302];\
        in_img_array[6][17][17] <= img[2303];\
        in_img_array[6][18][0] <= img[2304];\
        in_img_array[6][18][1] <= img[2305];\
        in_img_array[6][18][2] <= img[2306];\
        in_img_array[6][18][3] <= img[2307];\
        in_img_array[6][18][4] <= img[2308];\
        in_img_array[6][18][5] <= img[2309];\
        in_img_array[6][18][6] <= img[2310];\
        in_img_array[6][18][7] <= img[2311];\
        in_img_array[6][18][8] <= img[2312];\
        in_img_array[6][18][9] <= img[2313];\
        in_img_array[6][18][10] <= img[2314];\
        in_img_array[6][18][11] <= img[2315];\
        in_img_array[6][18][12] <= img[2316];\
        in_img_array[6][18][13] <= img[2317];\
        in_img_array[6][18][14] <= img[2318];\
        in_img_array[6][18][15] <= img[2319];\
        in_img_array[6][18][16] <= img[2320];\
        in_img_array[6][18][17] <= img[2321];\
        in_img_array[6][19][0] <= img[2322];\
        in_img_array[6][19][1] <= img[2323];\
        in_img_array[6][19][2] <= img[2324];\
        in_img_array[6][19][3] <= img[2325];\
        in_img_array[6][19][4] <= img[2326];\
        in_img_array[6][19][5] <= img[2327];\
        in_img_array[6][19][6] <= img[2328];\
        in_img_array[6][19][7] <= img[2329];\
        in_img_array[6][19][8] <= img[2330];\
        in_img_array[6][19][9] <= img[2331];\
        in_img_array[6][19][10] <= img[2332];\
        in_img_array[6][19][11] <= img[2333];\
        in_img_array[6][19][12] <= img[2334];\
        in_img_array[6][19][13] <= img[2335];\
        in_img_array[6][19][14] <= img[2336];\
        in_img_array[6][19][15] <= img[2337];\
        in_img_array[6][19][16] <= img[2338];\
        in_img_array[6][19][17] <= img[2339];\
        in_img_array[6][20][0] <= img[2340];\
        in_img_array[6][20][1] <= img[2341];\
        in_img_array[6][20][2] <= img[2342];\
        in_img_array[6][20][3] <= img[2343];\
        in_img_array[6][20][4] <= img[2344];\
        in_img_array[6][20][5] <= img[2345];\
        in_img_array[6][20][6] <= img[2346];\
        in_img_array[6][20][7] <= img[2347];\
        in_img_array[6][20][8] <= img[2348];\
        in_img_array[6][20][9] <= img[2349];\
        in_img_array[6][20][10] <= img[2350];\
        in_img_array[6][20][11] <= img[2351];\
        in_img_array[6][20][12] <= img[2352];\
        in_img_array[6][20][13] <= img[2353];\
        in_img_array[6][20][14] <= img[2354];\
        in_img_array[6][20][15] <= img[2355];\
        in_img_array[6][20][16] <= img[2356];\
        in_img_array[6][20][17] <= img[2357];\
        in_img_array[6][21][0] <= img[2358];\
        in_img_array[6][21][1] <= img[2359];\
        in_img_array[6][21][2] <= img[2360];\
        in_img_array[6][21][3] <= img[2361];\
        in_img_array[6][21][4] <= img[2362];\
        in_img_array[6][21][5] <= img[2363];\
        in_img_array[6][21][6] <= img[2364];\
        in_img_array[6][21][7] <= img[2365];\
        in_img_array[6][21][8] <= img[2366];\
        in_img_array[6][21][9] <= img[2367];\
        in_img_array[6][21][10] <= img[2368];\
        in_img_array[6][21][11] <= img[2369];\
        in_img_array[6][21][12] <= img[2370];\
        in_img_array[6][21][13] <= img[2371];\
        in_img_array[6][21][14] <= img[2372];\
        in_img_array[6][21][15] <= img[2373];\
        in_img_array[6][21][16] <= img[2374];\
        in_img_array[6][21][17] <= img[2375];\
        in_img_array[6][22][0] <= img[2376];\
        in_img_array[6][22][1] <= img[2377];\
        in_img_array[6][22][2] <= img[2378];\
        in_img_array[6][22][3] <= img[2379];\
        in_img_array[6][22][4] <= img[2380];\
        in_img_array[6][22][5] <= img[2381];\
        in_img_array[6][22][6] <= img[2382];\
        in_img_array[6][22][7] <= img[2383];\
        in_img_array[6][22][8] <= img[2384];\
        in_img_array[6][22][9] <= img[2385];\
        in_img_array[6][22][10] <= img[2386];\
        in_img_array[6][22][11] <= img[2387];\
        in_img_array[6][22][12] <= img[2388];\
        in_img_array[6][22][13] <= img[2389];\
        in_img_array[6][22][14] <= img[2390];\
        in_img_array[6][22][15] <= img[2391];\
        in_img_array[6][22][16] <= img[2392];\
        in_img_array[6][22][17] <= img[2393];\
        in_img_array[6][23][0] <= img[2394];\
        in_img_array[6][23][1] <= img[2395];\
        in_img_array[6][23][2] <= img[2396];\
        in_img_array[6][23][3] <= img[2397];\
        in_img_array[6][23][4] <= img[2398];\
        in_img_array[6][23][5] <= img[2399];\
        in_img_array[6][23][6] <= img[2400];\
        in_img_array[6][23][7] <= img[2401];\
        in_img_array[6][23][8] <= img[2402];\
        in_img_array[6][23][9] <= img[2403];\
        in_img_array[6][23][10] <= img[2404];\
        in_img_array[6][23][11] <= img[2405];\
        in_img_array[6][23][12] <= img[2406];\
        in_img_array[6][23][13] <= img[2407];\
        in_img_array[6][23][14] <= img[2408];\
        in_img_array[6][23][15] <= img[2409];\
        in_img_array[6][23][16] <= img[2410];\
        in_img_array[6][23][17] <= img[2411];\
        in_img_array[6][24][0] <= img[2412];\
        in_img_array[6][24][1] <= img[2413];\
        in_img_array[6][24][2] <= img[2414];\
        in_img_array[6][24][3] <= img[2415];\
        in_img_array[6][24][4] <= img[2416];\
        in_img_array[6][24][5] <= img[2417];\
        in_img_array[6][24][6] <= img[2418];\
        in_img_array[6][24][7] <= img[2419];\
        in_img_array[6][24][8] <= img[2420];\
        in_img_array[6][24][9] <= img[2421];\
        in_img_array[6][24][10] <= img[2422];\
        in_img_array[6][24][11] <= img[2423];\
        in_img_array[6][24][12] <= img[2424];\
        in_img_array[6][24][13] <= img[2425];\
        in_img_array[6][24][14] <= img[2426];\
        in_img_array[6][24][15] <= img[2427];\
        in_img_array[6][24][16] <= img[2428];\
        in_img_array[6][24][17] <= img[2429];\
        in_img_array[6][25][0] <= img[2430];\
        in_img_array[6][25][1] <= img[2431];\
        in_img_array[6][25][2] <= img[2432];\
        in_img_array[6][25][3] <= img[2433];\
        in_img_array[6][25][4] <= img[2434];\
        in_img_array[6][25][5] <= img[2435];\
        in_img_array[6][25][6] <= img[2436];\
        in_img_array[6][25][7] <= img[2437];\
        in_img_array[6][25][8] <= img[2438];\
        in_img_array[6][25][9] <= img[2439];\
        in_img_array[6][25][10] <= img[2440];\
        in_img_array[6][25][11] <= img[2441];\
        in_img_array[6][25][12] <= img[2442];\
        in_img_array[6][25][13] <= img[2443];\
        in_img_array[6][25][14] <= img[2444];\
        in_img_array[6][25][15] <= img[2445];\
        in_img_array[6][25][16] <= img[2446];\
        in_img_array[6][25][17] <= img[2447];\
        in_img_array[6][26][0] <= img[2448];\
        in_img_array[6][26][1] <= img[2449];\
        in_img_array[6][26][2] <= img[2450];\
        in_img_array[6][26][3] <= img[2451];\
        in_img_array[6][26][4] <= img[2452];\
        in_img_array[6][26][5] <= img[2453];\
        in_img_array[6][26][6] <= img[2454];\
        in_img_array[6][26][7] <= img[2455];\
        in_img_array[6][26][8] <= img[2456];\
        in_img_array[6][26][9] <= img[2457];\
        in_img_array[6][26][10] <= img[2458];\
        in_img_array[6][26][11] <= img[2459];\
        in_img_array[6][26][12] <= img[2460];\
        in_img_array[6][26][13] <= img[2461];\
        in_img_array[6][26][14] <= img[2462];\
        in_img_array[6][26][15] <= img[2463];\
        in_img_array[6][26][16] <= img[2464];\
        in_img_array[6][26][17] <= img[2465];\
        in_img_array[6][27][0] <= img[2466];\
        in_img_array[6][27][1] <= img[2467];\
        in_img_array[6][27][2] <= img[2468];\
        in_img_array[6][27][3] <= img[2469];\
        in_img_array[6][27][4] <= img[2470];\
        in_img_array[6][27][5] <= img[2471];\
        in_img_array[6][27][6] <= img[2472];\
        in_img_array[6][27][7] <= img[2473];\
        in_img_array[6][27][8] <= img[2474];\
        in_img_array[6][27][9] <= img[2475];\
        in_img_array[6][27][10] <= img[2476];\
        in_img_array[6][27][11] <= img[2477];\
        in_img_array[6][27][12] <= img[2478];\
        in_img_array[6][27][13] <= img[2479];\
        in_img_array[6][27][14] <= img[2480];\
        in_img_array[6][27][15] <= img[2481];\
        in_img_array[6][27][16] <= img[2482];\
        in_img_array[6][27][17] <= img[2483];\
        in_img_array[6][28][0] <= img[2484];\
        in_img_array[6][28][1] <= img[2485];\
        in_img_array[6][28][2] <= img[2486];\
        in_img_array[6][28][3] <= img[2487];\
        in_img_array[6][28][4] <= img[2488];\
        in_img_array[6][28][5] <= img[2489];\
        in_img_array[6][28][6] <= img[2490];\
        in_img_array[6][28][7] <= img[2491];\
        in_img_array[6][28][8] <= img[2492];\
        in_img_array[6][28][9] <= img[2493];\
        in_img_array[6][28][10] <= img[2494];\
        in_img_array[6][28][11] <= img[2495];\
        in_img_array[6][28][12] <= img[2496];\
        in_img_array[6][28][13] <= img[2497];\
        in_img_array[6][28][14] <= img[2498];\
        in_img_array[6][28][15] <= img[2499];\
        in_img_array[6][28][16] <= img[2500];\
        in_img_array[6][28][17] <= img[2501];\
        in_img_array[6][29][0] <= img[2502];\
        in_img_array[6][29][1] <= img[2503];\
        in_img_array[6][29][2] <= img[2504];\
        in_img_array[6][29][3] <= img[2505];\
        in_img_array[6][29][4] <= img[2506];\
        in_img_array[6][29][5] <= img[2507];\
        in_img_array[6][29][6] <= img[2508];\
        in_img_array[6][29][7] <= img[2509];\
        in_img_array[6][29][8] <= img[2510];\
        in_img_array[6][29][9] <= img[2511];\
        in_img_array[6][29][10] <= img[2512];\
        in_img_array[6][29][11] <= img[2513];\
        in_img_array[6][29][12] <= img[2514];\
        in_img_array[6][29][13] <= img[2515];\
        in_img_array[6][29][14] <= img[2516];\
        in_img_array[6][29][15] <= img[2517];\
        in_img_array[6][29][16] <= img[2518];\
        in_img_array[6][29][17] <= img[2519];\
        in_img_array[7][2][0] <= img[2520];\
        in_img_array[7][2][1] <= img[2521];\
        in_img_array[7][2][2] <= img[2522];\
        in_img_array[7][2][3] <= img[2523];\
        in_img_array[7][2][4] <= img[2524];\
        in_img_array[7][2][5] <= img[2525];\
        in_img_array[7][2][6] <= img[2526];\
        in_img_array[7][2][7] <= img[2527];\
        in_img_array[7][2][8] <= img[2528];\
        in_img_array[7][2][9] <= img[2529];\
        in_img_array[7][2][10] <= img[2530];\
        in_img_array[7][2][11] <= img[2531];\
        in_img_array[7][2][12] <= img[2532];\
        in_img_array[7][2][13] <= img[2533];\
        in_img_array[7][2][14] <= img[2534];\
        in_img_array[7][2][15] <= img[2535];\
        in_img_array[7][2][16] <= img[2536];\
        in_img_array[7][2][17] <= img[2537];\
        in_img_array[7][3][0] <= img[2538];\
        in_img_array[7][3][1] <= img[2539];\
        in_img_array[7][3][2] <= img[2540];\
        in_img_array[7][3][3] <= img[2541];\
        in_img_array[7][3][4] <= img[2542];\
        in_img_array[7][3][5] <= img[2543];\
        in_img_array[7][3][6] <= img[2544];\
        in_img_array[7][3][7] <= img[2545];\
        in_img_array[7][3][8] <= img[2546];\
        in_img_array[7][3][9] <= img[2547];\
        in_img_array[7][3][10] <= img[2548];\
        in_img_array[7][3][11] <= img[2549];\
        in_img_array[7][3][12] <= img[2550];\
        in_img_array[7][3][13] <= img[2551];\
        in_img_array[7][3][14] <= img[2552];\
        in_img_array[7][3][15] <= img[2553];\
        in_img_array[7][3][16] <= img[2554];\
        in_img_array[7][3][17] <= img[2555];\
        in_img_array[7][4][0] <= img[2556];\
        in_img_array[7][4][1] <= img[2557];\
        in_img_array[7][4][2] <= img[2558];\
        in_img_array[7][4][3] <= img[2559];\
        in_img_array[7][4][4] <= img[2560];\
        in_img_array[7][4][5] <= img[2561];\
        in_img_array[7][4][6] <= img[2562];\
        in_img_array[7][4][7] <= img[2563];\
        in_img_array[7][4][8] <= img[2564];\
        in_img_array[7][4][9] <= img[2565];\
        in_img_array[7][4][10] <= img[2566];\
        in_img_array[7][4][11] <= img[2567];\
        in_img_array[7][4][12] <= img[2568];\
        in_img_array[7][4][13] <= img[2569];\
        in_img_array[7][4][14] <= img[2570];\
        in_img_array[7][4][15] <= img[2571];\
        in_img_array[7][4][16] <= img[2572];\
        in_img_array[7][4][17] <= img[2573];\
        in_img_array[7][5][0] <= img[2574];\
        in_img_array[7][5][1] <= img[2575];\
        in_img_array[7][5][2] <= img[2576];\
        in_img_array[7][5][3] <= img[2577];\
        in_img_array[7][5][4] <= img[2578];\
        in_img_array[7][5][5] <= img[2579];\
        in_img_array[7][5][6] <= img[2580];\
        in_img_array[7][5][7] <= img[2581];\
        in_img_array[7][5][8] <= img[2582];\
        in_img_array[7][5][9] <= img[2583];\
        in_img_array[7][5][10] <= img[2584];\
        in_img_array[7][5][11] <= img[2585];\
        in_img_array[7][5][12] <= img[2586];\
        in_img_array[7][5][13] <= img[2587];\
        in_img_array[7][5][14] <= img[2588];\
        in_img_array[7][5][15] <= img[2589];\
        in_img_array[7][5][16] <= img[2590];\
        in_img_array[7][5][17] <= img[2591];\
        in_img_array[7][6][0] <= img[2592];\
        in_img_array[7][6][1] <= img[2593];\
        in_img_array[7][6][2] <= img[2594];\
        in_img_array[7][6][3] <= img[2595];\
        in_img_array[7][6][4] <= img[2596];\
        in_img_array[7][6][5] <= img[2597];\
        in_img_array[7][6][6] <= img[2598];\
        in_img_array[7][6][7] <= img[2599];\
        in_img_array[7][6][8] <= img[2600];\
        in_img_array[7][6][9] <= img[2601];\
        in_img_array[7][6][10] <= img[2602];\
        in_img_array[7][6][11] <= img[2603];\
        in_img_array[7][6][12] <= img[2604];\
        in_img_array[7][6][13] <= img[2605];\
        in_img_array[7][6][14] <= img[2606];\
        in_img_array[7][6][15] <= img[2607];\
        in_img_array[7][6][16] <= img[2608];\
        in_img_array[7][6][17] <= img[2609];\
        in_img_array[7][7][0] <= img[2610];\
        in_img_array[7][7][1] <= img[2611];\
        in_img_array[7][7][2] <= img[2612];\
        in_img_array[7][7][3] <= img[2613];\
        in_img_array[7][7][4] <= img[2614];\
        in_img_array[7][7][5] <= img[2615];\
        in_img_array[7][7][6] <= img[2616];\
        in_img_array[7][7][7] <= img[2617];\
        in_img_array[7][7][8] <= img[2618];\
        in_img_array[7][7][9] <= img[2619];\
        in_img_array[7][7][10] <= img[2620];\
        in_img_array[7][7][11] <= img[2621];\
        in_img_array[7][7][12] <= img[2622];\
        in_img_array[7][7][13] <= img[2623];\
        in_img_array[7][7][14] <= img[2624];\
        in_img_array[7][7][15] <= img[2625];\
        in_img_array[7][7][16] <= img[2626];\
        in_img_array[7][7][17] <= img[2627];\
        in_img_array[7][8][0] <= img[2628];\
        in_img_array[7][8][1] <= img[2629];\
        in_img_array[7][8][2] <= img[2630];\
        in_img_array[7][8][3] <= img[2631];\
        in_img_array[7][8][4] <= img[2632];\
        in_img_array[7][8][5] <= img[2633];\
        in_img_array[7][8][6] <= img[2634];\
        in_img_array[7][8][7] <= img[2635];\
        in_img_array[7][8][8] <= img[2636];\
        in_img_array[7][8][9] <= img[2637];\
        in_img_array[7][8][10] <= img[2638];\
        in_img_array[7][8][11] <= img[2639];\
        in_img_array[7][8][12] <= img[2640];\
        in_img_array[7][8][13] <= img[2641];\
        in_img_array[7][8][14] <= img[2642];\
        in_img_array[7][8][15] <= img[2643];\
        in_img_array[7][8][16] <= img[2644];\
        in_img_array[7][8][17] <= img[2645];\
        in_img_array[7][9][0] <= img[2646];\
        in_img_array[7][9][1] <= img[2647];\
        in_img_array[7][9][2] <= img[2648];\
        in_img_array[7][9][3] <= img[2649];\
        in_img_array[7][9][4] <= img[2650];\
        in_img_array[7][9][5] <= img[2651];\
        in_img_array[7][9][6] <= img[2652];\
        in_img_array[7][9][7] <= img[2653];\
        in_img_array[7][9][8] <= img[2654];\
        in_img_array[7][9][9] <= img[2655];\
        in_img_array[7][9][10] <= img[2656];\
        in_img_array[7][9][11] <= img[2657];\
        in_img_array[7][9][12] <= img[2658];\
        in_img_array[7][9][13] <= img[2659];\
        in_img_array[7][9][14] <= img[2660];\
        in_img_array[7][9][15] <= img[2661];\
        in_img_array[7][9][16] <= img[2662];\
        in_img_array[7][9][17] <= img[2663];\
        in_img_array[7][10][0] <= img[2664];\
        in_img_array[7][10][1] <= img[2665];\
        in_img_array[7][10][2] <= img[2666];\
        in_img_array[7][10][3] <= img[2667];\
        in_img_array[7][10][4] <= img[2668];\
        in_img_array[7][10][5] <= img[2669];\
        in_img_array[7][10][6] <= img[2670];\
        in_img_array[7][10][7] <= img[2671];\
        in_img_array[7][10][8] <= img[2672];\
        in_img_array[7][10][9] <= img[2673];\
        in_img_array[7][10][10] <= img[2674];\
        in_img_array[7][10][11] <= img[2675];\
        in_img_array[7][10][12] <= img[2676];\
        in_img_array[7][10][13] <= img[2677];\
        in_img_array[7][10][14] <= img[2678];\
        in_img_array[7][10][15] <= img[2679];\
        in_img_array[7][10][16] <= img[2680];\
        in_img_array[7][10][17] <= img[2681];\
        in_img_array[7][11][0] <= img[2682];\
        in_img_array[7][11][1] <= img[2683];\
        in_img_array[7][11][2] <= img[2684];\
        in_img_array[7][11][3] <= img[2685];\
        in_img_array[7][11][4] <= img[2686];\
        in_img_array[7][11][5] <= img[2687];\
        in_img_array[7][11][6] <= img[2688];\
        in_img_array[7][11][7] <= img[2689];\
        in_img_array[7][11][8] <= img[2690];\
        in_img_array[7][11][9] <= img[2691];\
        in_img_array[7][11][10] <= img[2692];\
        in_img_array[7][11][11] <= img[2693];\
        in_img_array[7][11][12] <= img[2694];\
        in_img_array[7][11][13] <= img[2695];\
        in_img_array[7][11][14] <= img[2696];\
        in_img_array[7][11][15] <= img[2697];\
        in_img_array[7][11][16] <= img[2698];\
        in_img_array[7][11][17] <= img[2699];\
        in_img_array[7][12][0] <= img[2700];\
        in_img_array[7][12][1] <= img[2701];\
        in_img_array[7][12][2] <= img[2702];\
        in_img_array[7][12][3] <= img[2703];\
        in_img_array[7][12][4] <= img[2704];\
        in_img_array[7][12][5] <= img[2705];\
        in_img_array[7][12][6] <= img[2706];\
        in_img_array[7][12][7] <= img[2707];\
        in_img_array[7][12][8] <= img[2708];\
        in_img_array[7][12][9] <= img[2709];\
        in_img_array[7][12][10] <= img[2710];\
        in_img_array[7][12][11] <= img[2711];\
        in_img_array[7][12][12] <= img[2712];\
        in_img_array[7][12][13] <= img[2713];\
        in_img_array[7][12][14] <= img[2714];\
        in_img_array[7][12][15] <= img[2715];\
        in_img_array[7][12][16] <= img[2716];\
        in_img_array[7][12][17] <= img[2717];\
        in_img_array[7][13][0] <= img[2718];\
        in_img_array[7][13][1] <= img[2719];\
        in_img_array[7][13][2] <= img[2720];\
        in_img_array[7][13][3] <= img[2721];\
        in_img_array[7][13][4] <= img[2722];\
        in_img_array[7][13][5] <= img[2723];\
        in_img_array[7][13][6] <= img[2724];\
        in_img_array[7][13][7] <= img[2725];\
        in_img_array[7][13][8] <= img[2726];\
        in_img_array[7][13][9] <= img[2727];\
        in_img_array[7][13][10] <= img[2728];\
        in_img_array[7][13][11] <= img[2729];\
        in_img_array[7][13][12] <= img[2730];\
        in_img_array[7][13][13] <= img[2731];\
        in_img_array[7][13][14] <= img[2732];\
        in_img_array[7][13][15] <= img[2733];\
        in_img_array[7][13][16] <= img[2734];\
        in_img_array[7][13][17] <= img[2735];\
        in_img_array[7][14][0] <= img[2736];\
        in_img_array[7][14][1] <= img[2737];\
        in_img_array[7][14][2] <= img[2738];\
        in_img_array[7][14][3] <= img[2739];\
        in_img_array[7][14][4] <= img[2740];\
        in_img_array[7][14][5] <= img[2741];\
        in_img_array[7][14][6] <= img[2742];\
        in_img_array[7][14][7] <= img[2743];\
        in_img_array[7][14][8] <= img[2744];\
        in_img_array[7][14][9] <= img[2745];\
        in_img_array[7][14][10] <= img[2746];\
        in_img_array[7][14][11] <= img[2747];\
        in_img_array[7][14][12] <= img[2748];\
        in_img_array[7][14][13] <= img[2749];\
        in_img_array[7][14][14] <= img[2750];\
        in_img_array[7][14][15] <= img[2751];\
        in_img_array[7][14][16] <= img[2752];\
        in_img_array[7][14][17] <= img[2753];\
        in_img_array[7][15][0] <= img[2754];\
        in_img_array[7][15][1] <= img[2755];\
        in_img_array[7][15][2] <= img[2756];\
        in_img_array[7][15][3] <= img[2757];\
        in_img_array[7][15][4] <= img[2758];\
        in_img_array[7][15][5] <= img[2759];\
        in_img_array[7][15][6] <= img[2760];\
        in_img_array[7][15][7] <= img[2761];\
        in_img_array[7][15][8] <= img[2762];\
        in_img_array[7][15][9] <= img[2763];\
        in_img_array[7][15][10] <= img[2764];\
        in_img_array[7][15][11] <= img[2765];\
        in_img_array[7][15][12] <= img[2766];\
        in_img_array[7][15][13] <= img[2767];\
        in_img_array[7][15][14] <= img[2768];\
        in_img_array[7][15][15] <= img[2769];\
        in_img_array[7][15][16] <= img[2770];\
        in_img_array[7][15][17] <= img[2771];\
        in_img_array[7][16][0] <= img[2772];\
        in_img_array[7][16][1] <= img[2773];\
        in_img_array[7][16][2] <= img[2774];\
        in_img_array[7][16][3] <= img[2775];\
        in_img_array[7][16][4] <= img[2776];\
        in_img_array[7][16][5] <= img[2777];\
        in_img_array[7][16][6] <= img[2778];\
        in_img_array[7][16][7] <= img[2779];\
        in_img_array[7][16][8] <= img[2780];\
        in_img_array[7][16][9] <= img[2781];\
        in_img_array[7][16][10] <= img[2782];\
        in_img_array[7][16][11] <= img[2783];\
        in_img_array[7][16][12] <= img[2784];\
        in_img_array[7][16][13] <= img[2785];\
        in_img_array[7][16][14] <= img[2786];\
        in_img_array[7][16][15] <= img[2787];\
        in_img_array[7][16][16] <= img[2788];\
        in_img_array[7][16][17] <= img[2789];\
        in_img_array[7][17][0] <= img[2790];\
        in_img_array[7][17][1] <= img[2791];\
        in_img_array[7][17][2] <= img[2792];\
        in_img_array[7][17][3] <= img[2793];\
        in_img_array[7][17][4] <= img[2794];\
        in_img_array[7][17][5] <= img[2795];\
        in_img_array[7][17][6] <= img[2796];\
        in_img_array[7][17][7] <= img[2797];\
        in_img_array[7][17][8] <= img[2798];\
        in_img_array[7][17][9] <= img[2799];\
        in_img_array[7][17][10] <= img[2800];\
        in_img_array[7][17][11] <= img[2801];\
        in_img_array[7][17][12] <= img[2802];\
        in_img_array[7][17][13] <= img[2803];\
        in_img_array[7][17][14] <= img[2804];\
        in_img_array[7][17][15] <= img[2805];\
        in_img_array[7][17][16] <= img[2806];\
        in_img_array[7][17][17] <= img[2807];\
        in_img_array[7][18][0] <= img[2808];\
        in_img_array[7][18][1] <= img[2809];\
        in_img_array[7][18][2] <= img[2810];\
        in_img_array[7][18][3] <= img[2811];\
        in_img_array[7][18][4] <= img[2812];\
        in_img_array[7][18][5] <= img[2813];\
        in_img_array[7][18][6] <= img[2814];\
        in_img_array[7][18][7] <= img[2815];\
        in_img_array[7][18][8] <= img[2816];\
        in_img_array[7][18][9] <= img[2817];\
        in_img_array[7][18][10] <= img[2818];\
        in_img_array[7][18][11] <= img[2819];\
        in_img_array[7][18][12] <= img[2820];\
        in_img_array[7][18][13] <= img[2821];\
        in_img_array[7][18][14] <= img[2822];\
        in_img_array[7][18][15] <= img[2823];\
        in_img_array[7][18][16] <= img[2824];\
        in_img_array[7][18][17] <= img[2825];\
        in_img_array[7][19][0] <= img[2826];\
        in_img_array[7][19][1] <= img[2827];\
        in_img_array[7][19][2] <= img[2828];\
        in_img_array[7][19][3] <= img[2829];\
        in_img_array[7][19][4] <= img[2830];\
        in_img_array[7][19][5] <= img[2831];\
        in_img_array[7][19][6] <= img[2832];\
        in_img_array[7][19][7] <= img[2833];\
        in_img_array[7][19][8] <= img[2834];\
        in_img_array[7][19][9] <= img[2835];\
        in_img_array[7][19][10] <= img[2836];\
        in_img_array[7][19][11] <= img[2837];\
        in_img_array[7][19][12] <= img[2838];\
        in_img_array[7][19][13] <= img[2839];\
        in_img_array[7][19][14] <= img[2840];\
        in_img_array[7][19][15] <= img[2841];\
        in_img_array[7][19][16] <= img[2842];\
        in_img_array[7][19][17] <= img[2843];\
        in_img_array[7][20][0] <= img[2844];\
        in_img_array[7][20][1] <= img[2845];\
        in_img_array[7][20][2] <= img[2846];\
        in_img_array[7][20][3] <= img[2847];\
        in_img_array[7][20][4] <= img[2848];\
        in_img_array[7][20][5] <= img[2849];\
        in_img_array[7][20][6] <= img[2850];\
        in_img_array[7][20][7] <= img[2851];\
        in_img_array[7][20][8] <= img[2852];\
        in_img_array[7][20][9] <= img[2853];\
        in_img_array[7][20][10] <= img[2854];\
        in_img_array[7][20][11] <= img[2855];\
        in_img_array[7][20][12] <= img[2856];\
        in_img_array[7][20][13] <= img[2857];\
        in_img_array[7][20][14] <= img[2858];\
        in_img_array[7][20][15] <= img[2859];\
        in_img_array[7][20][16] <= img[2860];\
        in_img_array[7][20][17] <= img[2861];\
        in_img_array[7][21][0] <= img[2862];\
        in_img_array[7][21][1] <= img[2863];\
        in_img_array[7][21][2] <= img[2864];\
        in_img_array[7][21][3] <= img[2865];\
        in_img_array[7][21][4] <= img[2866];\
        in_img_array[7][21][5] <= img[2867];\
        in_img_array[7][21][6] <= img[2868];\
        in_img_array[7][21][7] <= img[2869];\
        in_img_array[7][21][8] <= img[2870];\
        in_img_array[7][21][9] <= img[2871];\
        in_img_array[7][21][10] <= img[2872];\
        in_img_array[7][21][11] <= img[2873];\
        in_img_array[7][21][12] <= img[2874];\
        in_img_array[7][21][13] <= img[2875];\
        in_img_array[7][21][14] <= img[2876];\
        in_img_array[7][21][15] <= img[2877];\
        in_img_array[7][21][16] <= img[2878];\
        in_img_array[7][21][17] <= img[2879];\
        in_img_array[7][22][0] <= img[2880];\
        in_img_array[7][22][1] <= img[2881];\
        in_img_array[7][22][2] <= img[2882];\
        in_img_array[7][22][3] <= img[2883];\
        in_img_array[7][22][4] <= img[2884];\
        in_img_array[7][22][5] <= img[2885];\
        in_img_array[7][22][6] <= img[2886];\
        in_img_array[7][22][7] <= img[2887];\
        in_img_array[7][22][8] <= img[2888];\
        in_img_array[7][22][9] <= img[2889];\
        in_img_array[7][22][10] <= img[2890];\
        in_img_array[7][22][11] <= img[2891];\
        in_img_array[7][22][12] <= img[2892];\
        in_img_array[7][22][13] <= img[2893];\
        in_img_array[7][22][14] <= img[2894];\
        in_img_array[7][22][15] <= img[2895];\
        in_img_array[7][22][16] <= img[2896];\
        in_img_array[7][22][17] <= img[2897];\
        in_img_array[7][23][0] <= img[2898];\
        in_img_array[7][23][1] <= img[2899];\
        in_img_array[7][23][2] <= img[2900];\
        in_img_array[7][23][3] <= img[2901];\
        in_img_array[7][23][4] <= img[2902];\
        in_img_array[7][23][5] <= img[2903];\
        in_img_array[7][23][6] <= img[2904];\
        in_img_array[7][23][7] <= img[2905];\
        in_img_array[7][23][8] <= img[2906];\
        in_img_array[7][23][9] <= img[2907];\
        in_img_array[7][23][10] <= img[2908];\
        in_img_array[7][23][11] <= img[2909];\
        in_img_array[7][23][12] <= img[2910];\
        in_img_array[7][23][13] <= img[2911];\
        in_img_array[7][23][14] <= img[2912];\
        in_img_array[7][23][15] <= img[2913];\
        in_img_array[7][23][16] <= img[2914];\
        in_img_array[7][23][17] <= img[2915];\
        in_img_array[7][24][0] <= img[2916];\
        in_img_array[7][24][1] <= img[2917];\
        in_img_array[7][24][2] <= img[2918];\
        in_img_array[7][24][3] <= img[2919];\
        in_img_array[7][24][4] <= img[2920];\
        in_img_array[7][24][5] <= img[2921];\
        in_img_array[7][24][6] <= img[2922];\
        in_img_array[7][24][7] <= img[2923];\
        in_img_array[7][24][8] <= img[2924];\
        in_img_array[7][24][9] <= img[2925];\
        in_img_array[7][24][10] <= img[2926];\
        in_img_array[7][24][11] <= img[2927];\
        in_img_array[7][24][12] <= img[2928];\
        in_img_array[7][24][13] <= img[2929];\
        in_img_array[7][24][14] <= img[2930];\
        in_img_array[7][24][15] <= img[2931];\
        in_img_array[7][24][16] <= img[2932];\
        in_img_array[7][24][17] <= img[2933];\
        in_img_array[7][25][0] <= img[2934];\
        in_img_array[7][25][1] <= img[2935];\
        in_img_array[7][25][2] <= img[2936];\
        in_img_array[7][25][3] <= img[2937];\
        in_img_array[7][25][4] <= img[2938];\
        in_img_array[7][25][5] <= img[2939];\
        in_img_array[7][25][6] <= img[2940];\
        in_img_array[7][25][7] <= img[2941];\
        in_img_array[7][25][8] <= img[2942];\
        in_img_array[7][25][9] <= img[2943];\
        in_img_array[7][25][10] <= img[2944];\
        in_img_array[7][25][11] <= img[2945];\
        in_img_array[7][25][12] <= img[2946];\
        in_img_array[7][25][13] <= img[2947];\
        in_img_array[7][25][14] <= img[2948];\
        in_img_array[7][25][15] <= img[2949];\
        in_img_array[7][25][16] <= img[2950];\
        in_img_array[7][25][17] <= img[2951];\
        in_img_array[7][26][0] <= img[2952];\
        in_img_array[7][26][1] <= img[2953];\
        in_img_array[7][26][2] <= img[2954];\
        in_img_array[7][26][3] <= img[2955];\
        in_img_array[7][26][4] <= img[2956];\
        in_img_array[7][26][5] <= img[2957];\
        in_img_array[7][26][6] <= img[2958];\
        in_img_array[7][26][7] <= img[2959];\
        in_img_array[7][26][8] <= img[2960];\
        in_img_array[7][26][9] <= img[2961];\
        in_img_array[7][26][10] <= img[2962];\
        in_img_array[7][26][11] <= img[2963];\
        in_img_array[7][26][12] <= img[2964];\
        in_img_array[7][26][13] <= img[2965];\
        in_img_array[7][26][14] <= img[2966];\
        in_img_array[7][26][15] <= img[2967];\
        in_img_array[7][26][16] <= img[2968];\
        in_img_array[7][26][17] <= img[2969];\
        in_img_array[7][27][0] <= img[2970];\
        in_img_array[7][27][1] <= img[2971];\
        in_img_array[7][27][2] <= img[2972];\
        in_img_array[7][27][3] <= img[2973];\
        in_img_array[7][27][4] <= img[2974];\
        in_img_array[7][27][5] <= img[2975];\
        in_img_array[7][27][6] <= img[2976];\
        in_img_array[7][27][7] <= img[2977];\
        in_img_array[7][27][8] <= img[2978];\
        in_img_array[7][27][9] <= img[2979];\
        in_img_array[7][27][10] <= img[2980];\
        in_img_array[7][27][11] <= img[2981];\
        in_img_array[7][27][12] <= img[2982];\
        in_img_array[7][27][13] <= img[2983];\
        in_img_array[7][27][14] <= img[2984];\
        in_img_array[7][27][15] <= img[2985];\
        in_img_array[7][27][16] <= img[2986];\
        in_img_array[7][27][17] <= img[2987];\
        in_img_array[7][28][0] <= img[2988];\
        in_img_array[7][28][1] <= img[2989];\
        in_img_array[7][28][2] <= img[2990];\
        in_img_array[7][28][3] <= img[2991];\
        in_img_array[7][28][4] <= img[2992];\
        in_img_array[7][28][5] <= img[2993];\
        in_img_array[7][28][6] <= img[2994];\
        in_img_array[7][28][7] <= img[2995];\
        in_img_array[7][28][8] <= img[2996];\
        in_img_array[7][28][9] <= img[2997];\
        in_img_array[7][28][10] <= img[2998];\
        in_img_array[7][28][11] <= img[2999];\
        in_img_array[7][28][12] <= img[3000];\
        in_img_array[7][28][13] <= img[3001];\
        in_img_array[7][28][14] <= img[3002];\
        in_img_array[7][28][15] <= img[3003];\
        in_img_array[7][28][16] <= img[3004];\
        in_img_array[7][28][17] <= img[3005];\
        in_img_array[7][29][0] <= img[3006];\
        in_img_array[7][29][1] <= img[3007];\
        in_img_array[7][29][2] <= img[3008];\
        in_img_array[7][29][3] <= img[3009];\
        in_img_array[7][29][4] <= img[3010];\
        in_img_array[7][29][5] <= img[3011];\
        in_img_array[7][29][6] <= img[3012];\
        in_img_array[7][29][7] <= img[3013];\
        in_img_array[7][29][8] <= img[3014];\
        in_img_array[7][29][9] <= img[3015];\
        in_img_array[7][29][10] <= img[3016];\
        in_img_array[7][29][11] <= img[3017];\
        in_img_array[7][29][12] <= img[3018];\
        in_img_array[7][29][13] <= img[3019];\
        in_img_array[7][29][14] <= img[3020];\
        in_img_array[7][29][15] <= img[3021];\
        in_img_array[7][29][16] <= img[3022];\
        in_img_array[7][29][17] <= img[3023];\
        in_img_array[8][2][0] <= img[3024];\
        in_img_array[8][2][1] <= img[3025];\
        in_img_array[8][2][2] <= img[3026];\
        in_img_array[8][2][3] <= img[3027];\
        in_img_array[8][2][4] <= img[3028];\
        in_img_array[8][2][5] <= img[3029];\
        in_img_array[8][2][6] <= img[3030];\
        in_img_array[8][2][7] <= img[3031];\
        in_img_array[8][2][8] <= img[3032];\
        in_img_array[8][2][9] <= img[3033];\
        in_img_array[8][2][10] <= img[3034];\
        in_img_array[8][2][11] <= img[3035];\
        in_img_array[8][2][12] <= img[3036];\
        in_img_array[8][2][13] <= img[3037];\
        in_img_array[8][2][14] <= img[3038];\
        in_img_array[8][2][15] <= img[3039];\
        in_img_array[8][2][16] <= img[3040];\
        in_img_array[8][2][17] <= img[3041];\
        in_img_array[8][3][0] <= img[3042];\
        in_img_array[8][3][1] <= img[3043];\
        in_img_array[8][3][2] <= img[3044];\
        in_img_array[8][3][3] <= img[3045];\
        in_img_array[8][3][4] <= img[3046];\
        in_img_array[8][3][5] <= img[3047];\
        in_img_array[8][3][6] <= img[3048];\
        in_img_array[8][3][7] <= img[3049];\
        in_img_array[8][3][8] <= img[3050];\
        in_img_array[8][3][9] <= img[3051];\
        in_img_array[8][3][10] <= img[3052];\
        in_img_array[8][3][11] <= img[3053];\
        in_img_array[8][3][12] <= img[3054];\
        in_img_array[8][3][13] <= img[3055];\
        in_img_array[8][3][14] <= img[3056];\
        in_img_array[8][3][15] <= img[3057];\
        in_img_array[8][3][16] <= img[3058];\
        in_img_array[8][3][17] <= img[3059];\
        in_img_array[8][4][0] <= img[3060];\
        in_img_array[8][4][1] <= img[3061];\
        in_img_array[8][4][2] <= img[3062];\
        in_img_array[8][4][3] <= img[3063];\
        in_img_array[8][4][4] <= img[3064];\
        in_img_array[8][4][5] <= img[3065];\
        in_img_array[8][4][6] <= img[3066];\
        in_img_array[8][4][7] <= img[3067];\
        in_img_array[8][4][8] <= img[3068];\
        in_img_array[8][4][9] <= img[3069];\
        in_img_array[8][4][10] <= img[3070];\
        in_img_array[8][4][11] <= img[3071];\
        in_img_array[8][4][12] <= img[3072];\
        in_img_array[8][4][13] <= img[3073];\
        in_img_array[8][4][14] <= img[3074];\
        in_img_array[8][4][15] <= img[3075];\
        in_img_array[8][4][16] <= img[3076];\
        in_img_array[8][4][17] <= img[3077];\
        in_img_array[8][5][0] <= img[3078];\
        in_img_array[8][5][1] <= img[3079];\
        in_img_array[8][5][2] <= img[3080];\
        in_img_array[8][5][3] <= img[3081];\
        in_img_array[8][5][4] <= img[3082];\
        in_img_array[8][5][5] <= img[3083];\
        in_img_array[8][5][6] <= img[3084];\
        in_img_array[8][5][7] <= img[3085];\
        in_img_array[8][5][8] <= img[3086];\
        in_img_array[8][5][9] <= img[3087];\
        in_img_array[8][5][10] <= img[3088];\
        in_img_array[8][5][11] <= img[3089];\
        in_img_array[8][5][12] <= img[3090];\
        in_img_array[8][5][13] <= img[3091];\
        in_img_array[8][5][14] <= img[3092];\
        in_img_array[8][5][15] <= img[3093];\
        in_img_array[8][5][16] <= img[3094];\
        in_img_array[8][5][17] <= img[3095];\
        in_img_array[8][6][0] <= img[3096];\
        in_img_array[8][6][1] <= img[3097];\
        in_img_array[8][6][2] <= img[3098];\
        in_img_array[8][6][3] <= img[3099];\
        in_img_array[8][6][4] <= img[3100];\
        in_img_array[8][6][5] <= img[3101];\
        in_img_array[8][6][6] <= img[3102];\
        in_img_array[8][6][7] <= img[3103];\
        in_img_array[8][6][8] <= img[3104];\
        in_img_array[8][6][9] <= img[3105];\
        in_img_array[8][6][10] <= img[3106];\
        in_img_array[8][6][11] <= img[3107];\
        in_img_array[8][6][12] <= img[3108];\
        in_img_array[8][6][13] <= img[3109];\
        in_img_array[8][6][14] <= img[3110];\
        in_img_array[8][6][15] <= img[3111];\
        in_img_array[8][6][16] <= img[3112];\
        in_img_array[8][6][17] <= img[3113];\
        in_img_array[8][7][0] <= img[3114];\
        in_img_array[8][7][1] <= img[3115];\
        in_img_array[8][7][2] <= img[3116];\
        in_img_array[8][7][3] <= img[3117];\
        in_img_array[8][7][4] <= img[3118];\
        in_img_array[8][7][5] <= img[3119];\
        in_img_array[8][7][6] <= img[3120];\
        in_img_array[8][7][7] <= img[3121];\
        in_img_array[8][7][8] <= img[3122];\
        in_img_array[8][7][9] <= img[3123];\
        in_img_array[8][7][10] <= img[3124];\
        in_img_array[8][7][11] <= img[3125];\
        in_img_array[8][7][12] <= img[3126];\
        in_img_array[8][7][13] <= img[3127];\
        in_img_array[8][7][14] <= img[3128];\
        in_img_array[8][7][15] <= img[3129];\
        in_img_array[8][7][16] <= img[3130];\
        in_img_array[8][7][17] <= img[3131];\
        in_img_array[8][8][0] <= img[3132];\
        in_img_array[8][8][1] <= img[3133];\
        in_img_array[8][8][2] <= img[3134];\
        in_img_array[8][8][3] <= img[3135];\
        in_img_array[8][8][4] <= img[3136];\
        in_img_array[8][8][5] <= img[3137];\
        in_img_array[8][8][6] <= img[3138];\
        in_img_array[8][8][7] <= img[3139];\
        in_img_array[8][8][8] <= img[3140];\
        in_img_array[8][8][9] <= img[3141];\
        in_img_array[8][8][10] <= img[3142];\
        in_img_array[8][8][11] <= img[3143];\
        in_img_array[8][8][12] <= img[3144];\
        in_img_array[8][8][13] <= img[3145];\
        in_img_array[8][8][14] <= img[3146];\
        in_img_array[8][8][15] <= img[3147];\
        in_img_array[8][8][16] <= img[3148];\
        in_img_array[8][8][17] <= img[3149];\
        in_img_array[8][9][0] <= img[3150];\
        in_img_array[8][9][1] <= img[3151];\
        in_img_array[8][9][2] <= img[3152];\
        in_img_array[8][9][3] <= img[3153];\
        in_img_array[8][9][4] <= img[3154];\
        in_img_array[8][9][5] <= img[3155];\
        in_img_array[8][9][6] <= img[3156];\
        in_img_array[8][9][7] <= img[3157];\
        in_img_array[8][9][8] <= img[3158];\
        in_img_array[8][9][9] <= img[3159];\
        in_img_array[8][9][10] <= img[3160];\
        in_img_array[8][9][11] <= img[3161];\
        in_img_array[8][9][12] <= img[3162];\
        in_img_array[8][9][13] <= img[3163];\
        in_img_array[8][9][14] <= img[3164];\
        in_img_array[8][9][15] <= img[3165];\
        in_img_array[8][9][16] <= img[3166];\
        in_img_array[8][9][17] <= img[3167];\
        in_img_array[8][10][0] <= img[3168];\
        in_img_array[8][10][1] <= img[3169];\
        in_img_array[8][10][2] <= img[3170];\
        in_img_array[8][10][3] <= img[3171];\
        in_img_array[8][10][4] <= img[3172];\
        in_img_array[8][10][5] <= img[3173];\
        in_img_array[8][10][6] <= img[3174];\
        in_img_array[8][10][7] <= img[3175];\
        in_img_array[8][10][8] <= img[3176];\
        in_img_array[8][10][9] <= img[3177];\
        in_img_array[8][10][10] <= img[3178];\
        in_img_array[8][10][11] <= img[3179];\
        in_img_array[8][10][12] <= img[3180];\
        in_img_array[8][10][13] <= img[3181];\
        in_img_array[8][10][14] <= img[3182];\
        in_img_array[8][10][15] <= img[3183];\
        in_img_array[8][10][16] <= img[3184];\
        in_img_array[8][10][17] <= img[3185];\
        in_img_array[8][11][0] <= img[3186];\
        in_img_array[8][11][1] <= img[3187];\
        in_img_array[8][11][2] <= img[3188];\
        in_img_array[8][11][3] <= img[3189];\
        in_img_array[8][11][4] <= img[3190];\
        in_img_array[8][11][5] <= img[3191];\
        in_img_array[8][11][6] <= img[3192];\
        in_img_array[8][11][7] <= img[3193];\
        in_img_array[8][11][8] <= img[3194];\
        in_img_array[8][11][9] <= img[3195];\
        in_img_array[8][11][10] <= img[3196];\
        in_img_array[8][11][11] <= img[3197];\
        in_img_array[8][11][12] <= img[3198];\
        in_img_array[8][11][13] <= img[3199];\
        in_img_array[8][11][14] <= img[3200];\
        in_img_array[8][11][15] <= img[3201];\
        in_img_array[8][11][16] <= img[3202];\
        in_img_array[8][11][17] <= img[3203];\
        in_img_array[8][12][0] <= img[3204];\
        in_img_array[8][12][1] <= img[3205];\
        in_img_array[8][12][2] <= img[3206];\
        in_img_array[8][12][3] <= img[3207];\
        in_img_array[8][12][4] <= img[3208];\
        in_img_array[8][12][5] <= img[3209];\
        in_img_array[8][12][6] <= img[3210];\
        in_img_array[8][12][7] <= img[3211];\
        in_img_array[8][12][8] <= img[3212];\
        in_img_array[8][12][9] <= img[3213];\
        in_img_array[8][12][10] <= img[3214];\
        in_img_array[8][12][11] <= img[3215];\
        in_img_array[8][12][12] <= img[3216];\
        in_img_array[8][12][13] <= img[3217];\
        in_img_array[8][12][14] <= img[3218];\
        in_img_array[8][12][15] <= img[3219];\
        in_img_array[8][12][16] <= img[3220];\
        in_img_array[8][12][17] <= img[3221];\
        in_img_array[8][13][0] <= img[3222];\
        in_img_array[8][13][1] <= img[3223];\
        in_img_array[8][13][2] <= img[3224];\
        in_img_array[8][13][3] <= img[3225];\
        in_img_array[8][13][4] <= img[3226];\
        in_img_array[8][13][5] <= img[3227];\
        in_img_array[8][13][6] <= img[3228];\
        in_img_array[8][13][7] <= img[3229];\
        in_img_array[8][13][8] <= img[3230];\
        in_img_array[8][13][9] <= img[3231];\
        in_img_array[8][13][10] <= img[3232];\
        in_img_array[8][13][11] <= img[3233];\
        in_img_array[8][13][12] <= img[3234];\
        in_img_array[8][13][13] <= img[3235];\
        in_img_array[8][13][14] <= img[3236];\
        in_img_array[8][13][15] <= img[3237];\
        in_img_array[8][13][16] <= img[3238];\
        in_img_array[8][13][17] <= img[3239];\
        in_img_array[8][14][0] <= img[3240];\
        in_img_array[8][14][1] <= img[3241];\
        in_img_array[8][14][2] <= img[3242];\
        in_img_array[8][14][3] <= img[3243];\
        in_img_array[8][14][4] <= img[3244];\
        in_img_array[8][14][5] <= img[3245];\
        in_img_array[8][14][6] <= img[3246];\
        in_img_array[8][14][7] <= img[3247];\
        in_img_array[8][14][8] <= img[3248];\
        in_img_array[8][14][9] <= img[3249];\
        in_img_array[8][14][10] <= img[3250];\
        in_img_array[8][14][11] <= img[3251];\
        in_img_array[8][14][12] <= img[3252];\
        in_img_array[8][14][13] <= img[3253];\
        in_img_array[8][14][14] <= img[3254];\
        in_img_array[8][14][15] <= img[3255];\
        in_img_array[8][14][16] <= img[3256];\
        in_img_array[8][14][17] <= img[3257];\
        in_img_array[8][15][0] <= img[3258];\
        in_img_array[8][15][1] <= img[3259];\
        in_img_array[8][15][2] <= img[3260];\
        in_img_array[8][15][3] <= img[3261];\
        in_img_array[8][15][4] <= img[3262];\
        in_img_array[8][15][5] <= img[3263];\
        in_img_array[8][15][6] <= img[3264];\
        in_img_array[8][15][7] <= img[3265];\
        in_img_array[8][15][8] <= img[3266];\
        in_img_array[8][15][9] <= img[3267];\
        in_img_array[8][15][10] <= img[3268];\
        in_img_array[8][15][11] <= img[3269];\
        in_img_array[8][15][12] <= img[3270];\
        in_img_array[8][15][13] <= img[3271];\
        in_img_array[8][15][14] <= img[3272];\
        in_img_array[8][15][15] <= img[3273];\
        in_img_array[8][15][16] <= img[3274];\
        in_img_array[8][15][17] <= img[3275];\
        in_img_array[8][16][0] <= img[3276];\
        in_img_array[8][16][1] <= img[3277];\
        in_img_array[8][16][2] <= img[3278];\
        in_img_array[8][16][3] <= img[3279];\
        in_img_array[8][16][4] <= img[3280];\
        in_img_array[8][16][5] <= img[3281];\
        in_img_array[8][16][6] <= img[3282];\
        in_img_array[8][16][7] <= img[3283];\
        in_img_array[8][16][8] <= img[3284];\
        in_img_array[8][16][9] <= img[3285];\
        in_img_array[8][16][10] <= img[3286];\
        in_img_array[8][16][11] <= img[3287];\
        in_img_array[8][16][12] <= img[3288];\
        in_img_array[8][16][13] <= img[3289];\
        in_img_array[8][16][14] <= img[3290];\
        in_img_array[8][16][15] <= img[3291];\
        in_img_array[8][16][16] <= img[3292];\
        in_img_array[8][16][17] <= img[3293];\
        in_img_array[8][17][0] <= img[3294];\
        in_img_array[8][17][1] <= img[3295];\
        in_img_array[8][17][2] <= img[3296];\
        in_img_array[8][17][3] <= img[3297];\
        in_img_array[8][17][4] <= img[3298];\
        in_img_array[8][17][5] <= img[3299];\
        in_img_array[8][17][6] <= img[3300];\
        in_img_array[8][17][7] <= img[3301];\
        in_img_array[8][17][8] <= img[3302];\
        in_img_array[8][17][9] <= img[3303];\
        in_img_array[8][17][10] <= img[3304];\
        in_img_array[8][17][11] <= img[3305];\
        in_img_array[8][17][12] <= img[3306];\
        in_img_array[8][17][13] <= img[3307];\
        in_img_array[8][17][14] <= img[3308];\
        in_img_array[8][17][15] <= img[3309];\
        in_img_array[8][17][16] <= img[3310];\
        in_img_array[8][17][17] <= img[3311];\
        in_img_array[8][18][0] <= img[3312];\
        in_img_array[8][18][1] <= img[3313];\
        in_img_array[8][18][2] <= img[3314];\
        in_img_array[8][18][3] <= img[3315];\
        in_img_array[8][18][4] <= img[3316];\
        in_img_array[8][18][5] <= img[3317];\
        in_img_array[8][18][6] <= img[3318];\
        in_img_array[8][18][7] <= img[3319];\
        in_img_array[8][18][8] <= img[3320];\
        in_img_array[8][18][9] <= img[3321];\
        in_img_array[8][18][10] <= img[3322];\
        in_img_array[8][18][11] <= img[3323];\
        in_img_array[8][18][12] <= img[3324];\
        in_img_array[8][18][13] <= img[3325];\
        in_img_array[8][18][14] <= img[3326];\
        in_img_array[8][18][15] <= img[3327];\
        in_img_array[8][18][16] <= img[3328];\
        in_img_array[8][18][17] <= img[3329];\
        in_img_array[8][19][0] <= img[3330];\
        in_img_array[8][19][1] <= img[3331];\
        in_img_array[8][19][2] <= img[3332];\
        in_img_array[8][19][3] <= img[3333];\
        in_img_array[8][19][4] <= img[3334];\
        in_img_array[8][19][5] <= img[3335];\
        in_img_array[8][19][6] <= img[3336];\
        in_img_array[8][19][7] <= img[3337];\
        in_img_array[8][19][8] <= img[3338];\
        in_img_array[8][19][9] <= img[3339];\
        in_img_array[8][19][10] <= img[3340];\
        in_img_array[8][19][11] <= img[3341];\
        in_img_array[8][19][12] <= img[3342];\
        in_img_array[8][19][13] <= img[3343];\
        in_img_array[8][19][14] <= img[3344];\
        in_img_array[8][19][15] <= img[3345];\
        in_img_array[8][19][16] <= img[3346];\
        in_img_array[8][19][17] <= img[3347];\
        in_img_array[8][20][0] <= img[3348];\
        in_img_array[8][20][1] <= img[3349];\
        in_img_array[8][20][2] <= img[3350];\
        in_img_array[8][20][3] <= img[3351];\
        in_img_array[8][20][4] <= img[3352];\
        in_img_array[8][20][5] <= img[3353];\
        in_img_array[8][20][6] <= img[3354];\
        in_img_array[8][20][7] <= img[3355];\
        in_img_array[8][20][8] <= img[3356];\
        in_img_array[8][20][9] <= img[3357];\
        in_img_array[8][20][10] <= img[3358];\
        in_img_array[8][20][11] <= img[3359];\
        in_img_array[8][20][12] <= img[3360];\
        in_img_array[8][20][13] <= img[3361];\
        in_img_array[8][20][14] <= img[3362];\
        in_img_array[8][20][15] <= img[3363];\
        in_img_array[8][20][16] <= img[3364];\
        in_img_array[8][20][17] <= img[3365];\
        in_img_array[8][21][0] <= img[3366];\
        in_img_array[8][21][1] <= img[3367];\
        in_img_array[8][21][2] <= img[3368];\
        in_img_array[8][21][3] <= img[3369];\
        in_img_array[8][21][4] <= img[3370];\
        in_img_array[8][21][5] <= img[3371];\
        in_img_array[8][21][6] <= img[3372];\
        in_img_array[8][21][7] <= img[3373];\
        in_img_array[8][21][8] <= img[3374];\
        in_img_array[8][21][9] <= img[3375];\
        in_img_array[8][21][10] <= img[3376];\
        in_img_array[8][21][11] <= img[3377];\
        in_img_array[8][21][12] <= img[3378];\
        in_img_array[8][21][13] <= img[3379];\
        in_img_array[8][21][14] <= img[3380];\
        in_img_array[8][21][15] <= img[3381];\
        in_img_array[8][21][16] <= img[3382];\
        in_img_array[8][21][17] <= img[3383];\
        in_img_array[8][22][0] <= img[3384];\
        in_img_array[8][22][1] <= img[3385];\
        in_img_array[8][22][2] <= img[3386];\
        in_img_array[8][22][3] <= img[3387];\
        in_img_array[8][22][4] <= img[3388];\
        in_img_array[8][22][5] <= img[3389];\
        in_img_array[8][22][6] <= img[3390];\
        in_img_array[8][22][7] <= img[3391];\
        in_img_array[8][22][8] <= img[3392];\
        in_img_array[8][22][9] <= img[3393];\
        in_img_array[8][22][10] <= img[3394];\
        in_img_array[8][22][11] <= img[3395];\
        in_img_array[8][22][12] <= img[3396];\
        in_img_array[8][22][13] <= img[3397];\
        in_img_array[8][22][14] <= img[3398];\
        in_img_array[8][22][15] <= img[3399];\
        in_img_array[8][22][16] <= img[3400];\
        in_img_array[8][22][17] <= img[3401];\
        in_img_array[8][23][0] <= img[3402];\
        in_img_array[8][23][1] <= img[3403];\
        in_img_array[8][23][2] <= img[3404];\
        in_img_array[8][23][3] <= img[3405];\
        in_img_array[8][23][4] <= img[3406];\
        in_img_array[8][23][5] <= img[3407];\
        in_img_array[8][23][6] <= img[3408];\
        in_img_array[8][23][7] <= img[3409];\
        in_img_array[8][23][8] <= img[3410];\
        in_img_array[8][23][9] <= img[3411];\
        in_img_array[8][23][10] <= img[3412];\
        in_img_array[8][23][11] <= img[3413];\
        in_img_array[8][23][12] <= img[3414];\
        in_img_array[8][23][13] <= img[3415];\
        in_img_array[8][23][14] <= img[3416];\
        in_img_array[8][23][15] <= img[3417];\
        in_img_array[8][23][16] <= img[3418];\
        in_img_array[8][23][17] <= img[3419];\
        in_img_array[8][24][0] <= img[3420];\
        in_img_array[8][24][1] <= img[3421];\
        in_img_array[8][24][2] <= img[3422];\
        in_img_array[8][24][3] <= img[3423];\
        in_img_array[8][24][4] <= img[3424];\
        in_img_array[8][24][5] <= img[3425];\
        in_img_array[8][24][6] <= img[3426];\
        in_img_array[8][24][7] <= img[3427];\
        in_img_array[8][24][8] <= img[3428];\
        in_img_array[8][24][9] <= img[3429];\
        in_img_array[8][24][10] <= img[3430];\
        in_img_array[8][24][11] <= img[3431];\
        in_img_array[8][24][12] <= img[3432];\
        in_img_array[8][24][13] <= img[3433];\
        in_img_array[8][24][14] <= img[3434];\
        in_img_array[8][24][15] <= img[3435];\
        in_img_array[8][24][16] <= img[3436];\
        in_img_array[8][24][17] <= img[3437];\
        in_img_array[8][25][0] <= img[3438];\
        in_img_array[8][25][1] <= img[3439];\
        in_img_array[8][25][2] <= img[3440];\
        in_img_array[8][25][3] <= img[3441];\
        in_img_array[8][25][4] <= img[3442];\
        in_img_array[8][25][5] <= img[3443];\
        in_img_array[8][25][6] <= img[3444];\
        in_img_array[8][25][7] <= img[3445];\
        in_img_array[8][25][8] <= img[3446];\
        in_img_array[8][25][9] <= img[3447];\
        in_img_array[8][25][10] <= img[3448];\
        in_img_array[8][25][11] <= img[3449];\
        in_img_array[8][25][12] <= img[3450];\
        in_img_array[8][25][13] <= img[3451];\
        in_img_array[8][25][14] <= img[3452];\
        in_img_array[8][25][15] <= img[3453];\
        in_img_array[8][25][16] <= img[3454];\
        in_img_array[8][25][17] <= img[3455];\
        in_img_array[8][26][0] <= img[3456];\
        in_img_array[8][26][1] <= img[3457];\
        in_img_array[8][26][2] <= img[3458];\
        in_img_array[8][26][3] <= img[3459];\
        in_img_array[8][26][4] <= img[3460];\
        in_img_array[8][26][5] <= img[3461];\
        in_img_array[8][26][6] <= img[3462];\
        in_img_array[8][26][7] <= img[3463];\
        in_img_array[8][26][8] <= img[3464];\
        in_img_array[8][26][9] <= img[3465];\
        in_img_array[8][26][10] <= img[3466];\
        in_img_array[8][26][11] <= img[3467];\
        in_img_array[8][26][12] <= img[3468];\
        in_img_array[8][26][13] <= img[3469];\
        in_img_array[8][26][14] <= img[3470];\
        in_img_array[8][26][15] <= img[3471];\
        in_img_array[8][26][16] <= img[3472];\
        in_img_array[8][26][17] <= img[3473];\
        in_img_array[8][27][0] <= img[3474];\
        in_img_array[8][27][1] <= img[3475];\
        in_img_array[8][27][2] <= img[3476];\
        in_img_array[8][27][3] <= img[3477];\
        in_img_array[8][27][4] <= img[3478];\
        in_img_array[8][27][5] <= img[3479];\
        in_img_array[8][27][6] <= img[3480];\
        in_img_array[8][27][7] <= img[3481];\
        in_img_array[8][27][8] <= img[3482];\
        in_img_array[8][27][9] <= img[3483];\
        in_img_array[8][27][10] <= img[3484];\
        in_img_array[8][27][11] <= img[3485];\
        in_img_array[8][27][12] <= img[3486];\
        in_img_array[8][27][13] <= img[3487];\
        in_img_array[8][27][14] <= img[3488];\
        in_img_array[8][27][15] <= img[3489];\
        in_img_array[8][27][16] <= img[3490];\
        in_img_array[8][27][17] <= img[3491];\
        in_img_array[8][28][0] <= img[3492];\
        in_img_array[8][28][1] <= img[3493];\
        in_img_array[8][28][2] <= img[3494];\
        in_img_array[8][28][3] <= img[3495];\
        in_img_array[8][28][4] <= img[3496];\
        in_img_array[8][28][5] <= img[3497];\
        in_img_array[8][28][6] <= img[3498];\
        in_img_array[8][28][7] <= img[3499];\
        in_img_array[8][28][8] <= img[3500];\
        in_img_array[8][28][9] <= img[3501];\
        in_img_array[8][28][10] <= img[3502];\
        in_img_array[8][28][11] <= img[3503];\
        in_img_array[8][28][12] <= img[3504];\
        in_img_array[8][28][13] <= img[3505];\
        in_img_array[8][28][14] <= img[3506];\
        in_img_array[8][28][15] <= img[3507];\
        in_img_array[8][28][16] <= img[3508];\
        in_img_array[8][28][17] <= img[3509];\
        in_img_array[8][29][0] <= img[3510];\
        in_img_array[8][29][1] <= img[3511];\
        in_img_array[8][29][2] <= img[3512];\
        in_img_array[8][29][3] <= img[3513];\
        in_img_array[8][29][4] <= img[3514];\
        in_img_array[8][29][5] <= img[3515];\
        in_img_array[8][29][6] <= img[3516];\
        in_img_array[8][29][7] <= img[3517];\
        in_img_array[8][29][8] <= img[3518];\
        in_img_array[8][29][9] <= img[3519];\
        in_img_array[8][29][10] <= img[3520];\
        in_img_array[8][29][11] <= img[3521];\
        in_img_array[8][29][12] <= img[3522];\
        in_img_array[8][29][13] <= img[3523];\
        in_img_array[8][29][14] <= img[3524];\
        in_img_array[8][29][15] <= img[3525];\
        in_img_array[8][29][16] <= img[3526];\
        in_img_array[8][29][17] <= img[3527];\
        in_img_array[9][2][0] <= img[3528];\
        in_img_array[9][2][1] <= img[3529];\
        in_img_array[9][2][2] <= img[3530];\
        in_img_array[9][2][3] <= img[3531];\
        in_img_array[9][2][4] <= img[3532];\
        in_img_array[9][2][5] <= img[3533];\
        in_img_array[9][2][6] <= img[3534];\
        in_img_array[9][2][7] <= img[3535];\
        in_img_array[9][2][8] <= img[3536];\
        in_img_array[9][2][9] <= img[3537];\
        in_img_array[9][2][10] <= img[3538];\
        in_img_array[9][2][11] <= img[3539];\
        in_img_array[9][2][12] <= img[3540];\
        in_img_array[9][2][13] <= img[3541];\
        in_img_array[9][2][14] <= img[3542];\
        in_img_array[9][2][15] <= img[3543];\
        in_img_array[9][2][16] <= img[3544];\
        in_img_array[9][2][17] <= img[3545];\
        in_img_array[9][3][0] <= img[3546];\
        in_img_array[9][3][1] <= img[3547];\
        in_img_array[9][3][2] <= img[3548];\
        in_img_array[9][3][3] <= img[3549];\
        in_img_array[9][3][4] <= img[3550];\
        in_img_array[9][3][5] <= img[3551];\
        in_img_array[9][3][6] <= img[3552];\
        in_img_array[9][3][7] <= img[3553];\
        in_img_array[9][3][8] <= img[3554];\
        in_img_array[9][3][9] <= img[3555];\
        in_img_array[9][3][10] <= img[3556];\
        in_img_array[9][3][11] <= img[3557];\
        in_img_array[9][3][12] <= img[3558];\
        in_img_array[9][3][13] <= img[3559];\
        in_img_array[9][3][14] <= img[3560];\
        in_img_array[9][3][15] <= img[3561];\
        in_img_array[9][3][16] <= img[3562];\
        in_img_array[9][3][17] <= img[3563];\
        in_img_array[9][4][0] <= img[3564];\
        in_img_array[9][4][1] <= img[3565];\
        in_img_array[9][4][2] <= img[3566];\
        in_img_array[9][4][3] <= img[3567];\
        in_img_array[9][4][4] <= img[3568];\
        in_img_array[9][4][5] <= img[3569];\
        in_img_array[9][4][6] <= img[3570];\
        in_img_array[9][4][7] <= img[3571];\
        in_img_array[9][4][8] <= img[3572];\
        in_img_array[9][4][9] <= img[3573];\
        in_img_array[9][4][10] <= img[3574];\
        in_img_array[9][4][11] <= img[3575];\
        in_img_array[9][4][12] <= img[3576];\
        in_img_array[9][4][13] <= img[3577];\
        in_img_array[9][4][14] <= img[3578];\
        in_img_array[9][4][15] <= img[3579];\
        in_img_array[9][4][16] <= img[3580];\
        in_img_array[9][4][17] <= img[3581];\
        in_img_array[9][5][0] <= img[3582];\
        in_img_array[9][5][1] <= img[3583];\
        in_img_array[9][5][2] <= img[3584];\
        in_img_array[9][5][3] <= img[3585];\
        in_img_array[9][5][4] <= img[3586];\
        in_img_array[9][5][5] <= img[3587];\
        in_img_array[9][5][6] <= img[3588];\
        in_img_array[9][5][7] <= img[3589];\
        in_img_array[9][5][8] <= img[3590];\
        in_img_array[9][5][9] <= img[3591];\
        in_img_array[9][5][10] <= img[3592];\
        in_img_array[9][5][11] <= img[3593];\
        in_img_array[9][5][12] <= img[3594];\
        in_img_array[9][5][13] <= img[3595];\
        in_img_array[9][5][14] <= img[3596];\
        in_img_array[9][5][15] <= img[3597];\
        in_img_array[9][5][16] <= img[3598];\
        in_img_array[9][5][17] <= img[3599];\
        in_img_array[9][6][0] <= img[3600];\
        in_img_array[9][6][1] <= img[3601];\
        in_img_array[9][6][2] <= img[3602];\
        in_img_array[9][6][3] <= img[3603];\
        in_img_array[9][6][4] <= img[3604];\
        in_img_array[9][6][5] <= img[3605];\
        in_img_array[9][6][6] <= img[3606];\
        in_img_array[9][6][7] <= img[3607];\
        in_img_array[9][6][8] <= img[3608];\
        in_img_array[9][6][9] <= img[3609];\
        in_img_array[9][6][10] <= img[3610];\
        in_img_array[9][6][11] <= img[3611];\
        in_img_array[9][6][12] <= img[3612];\
        in_img_array[9][6][13] <= img[3613];\
        in_img_array[9][6][14] <= img[3614];\
        in_img_array[9][6][15] <= img[3615];\
        in_img_array[9][6][16] <= img[3616];\
        in_img_array[9][6][17] <= img[3617];\
        in_img_array[9][7][0] <= img[3618];\
        in_img_array[9][7][1] <= img[3619];\
        in_img_array[9][7][2] <= img[3620];\
        in_img_array[9][7][3] <= img[3621];\
        in_img_array[9][7][4] <= img[3622];\
        in_img_array[9][7][5] <= img[3623];\
        in_img_array[9][7][6] <= img[3624];\
        in_img_array[9][7][7] <= img[3625];\
        in_img_array[9][7][8] <= img[3626];\
        in_img_array[9][7][9] <= img[3627];\
        in_img_array[9][7][10] <= img[3628];\
        in_img_array[9][7][11] <= img[3629];\
        in_img_array[9][7][12] <= img[3630];\
        in_img_array[9][7][13] <= img[3631];\
        in_img_array[9][7][14] <= img[3632];\
        in_img_array[9][7][15] <= img[3633];\
        in_img_array[9][7][16] <= img[3634];\
        in_img_array[9][7][17] <= img[3635];\
        in_img_array[9][8][0] <= img[3636];\
        in_img_array[9][8][1] <= img[3637];\
        in_img_array[9][8][2] <= img[3638];\
        in_img_array[9][8][3] <= img[3639];\
        in_img_array[9][8][4] <= img[3640];\
        in_img_array[9][8][5] <= img[3641];\
        in_img_array[9][8][6] <= img[3642];\
        in_img_array[9][8][7] <= img[3643];\
        in_img_array[9][8][8] <= img[3644];\
        in_img_array[9][8][9] <= img[3645];\
        in_img_array[9][8][10] <= img[3646];\
        in_img_array[9][8][11] <= img[3647];\
        in_img_array[9][8][12] <= img[3648];\
        in_img_array[9][8][13] <= img[3649];\
        in_img_array[9][8][14] <= img[3650];\
        in_img_array[9][8][15] <= img[3651];\
        in_img_array[9][8][16] <= img[3652];\
        in_img_array[9][8][17] <= img[3653];\
        in_img_array[9][9][0] <= img[3654];\
        in_img_array[9][9][1] <= img[3655];\
        in_img_array[9][9][2] <= img[3656];\
        in_img_array[9][9][3] <= img[3657];\
        in_img_array[9][9][4] <= img[3658];\
        in_img_array[9][9][5] <= img[3659];\
        in_img_array[9][9][6] <= img[3660];\
        in_img_array[9][9][7] <= img[3661];\
        in_img_array[9][9][8] <= img[3662];\
        in_img_array[9][9][9] <= img[3663];\
        in_img_array[9][9][10] <= img[3664];\
        in_img_array[9][9][11] <= img[3665];\
        in_img_array[9][9][12] <= img[3666];\
        in_img_array[9][9][13] <= img[3667];\
        in_img_array[9][9][14] <= img[3668];\
        in_img_array[9][9][15] <= img[3669];\
        in_img_array[9][9][16] <= img[3670];\
        in_img_array[9][9][17] <= img[3671];\
        in_img_array[9][10][0] <= img[3672];\
        in_img_array[9][10][1] <= img[3673];\
        in_img_array[9][10][2] <= img[3674];\
        in_img_array[9][10][3] <= img[3675];\
        in_img_array[9][10][4] <= img[3676];\
        in_img_array[9][10][5] <= img[3677];\
        in_img_array[9][10][6] <= img[3678];\
        in_img_array[9][10][7] <= img[3679];\
        in_img_array[9][10][8] <= img[3680];\
        in_img_array[9][10][9] <= img[3681];\
        in_img_array[9][10][10] <= img[3682];\
        in_img_array[9][10][11] <= img[3683];\
        in_img_array[9][10][12] <= img[3684];\
        in_img_array[9][10][13] <= img[3685];\
        in_img_array[9][10][14] <= img[3686];\
        in_img_array[9][10][15] <= img[3687];\
        in_img_array[9][10][16] <= img[3688];\
        in_img_array[9][10][17] <= img[3689];\
        in_img_array[9][11][0] <= img[3690];\
        in_img_array[9][11][1] <= img[3691];\
        in_img_array[9][11][2] <= img[3692];\
        in_img_array[9][11][3] <= img[3693];\
        in_img_array[9][11][4] <= img[3694];\
        in_img_array[9][11][5] <= img[3695];\
        in_img_array[9][11][6] <= img[3696];\
        in_img_array[9][11][7] <= img[3697];\
        in_img_array[9][11][8] <= img[3698];\
        in_img_array[9][11][9] <= img[3699];\
        in_img_array[9][11][10] <= img[3700];\
        in_img_array[9][11][11] <= img[3701];\
        in_img_array[9][11][12] <= img[3702];\
        in_img_array[9][11][13] <= img[3703];\
        in_img_array[9][11][14] <= img[3704];\
        in_img_array[9][11][15] <= img[3705];\
        in_img_array[9][11][16] <= img[3706];\
        in_img_array[9][11][17] <= img[3707];\
        in_img_array[9][12][0] <= img[3708];\
        in_img_array[9][12][1] <= img[3709];\
        in_img_array[9][12][2] <= img[3710];\
        in_img_array[9][12][3] <= img[3711];\
        in_img_array[9][12][4] <= img[3712];\
        in_img_array[9][12][5] <= img[3713];\
        in_img_array[9][12][6] <= img[3714];\
        in_img_array[9][12][7] <= img[3715];\
        in_img_array[9][12][8] <= img[3716];\
        in_img_array[9][12][9] <= img[3717];\
        in_img_array[9][12][10] <= img[3718];\
        in_img_array[9][12][11] <= img[3719];\
        in_img_array[9][12][12] <= img[3720];\
        in_img_array[9][12][13] <= img[3721];\
        in_img_array[9][12][14] <= img[3722];\
        in_img_array[9][12][15] <= img[3723];\
        in_img_array[9][12][16] <= img[3724];\
        in_img_array[9][12][17] <= img[3725];\
        in_img_array[9][13][0] <= img[3726];\
        in_img_array[9][13][1] <= img[3727];\
        in_img_array[9][13][2] <= img[3728];\
        in_img_array[9][13][3] <= img[3729];\
        in_img_array[9][13][4] <= img[3730];\
        in_img_array[9][13][5] <= img[3731];\
        in_img_array[9][13][6] <= img[3732];\
        in_img_array[9][13][7] <= img[3733];\
        in_img_array[9][13][8] <= img[3734];\
        in_img_array[9][13][9] <= img[3735];\
        in_img_array[9][13][10] <= img[3736];\
        in_img_array[9][13][11] <= img[3737];\
        in_img_array[9][13][12] <= img[3738];\
        in_img_array[9][13][13] <= img[3739];\
        in_img_array[9][13][14] <= img[3740];\
        in_img_array[9][13][15] <= img[3741];\
        in_img_array[9][13][16] <= img[3742];\
        in_img_array[9][13][17] <= img[3743];\
        in_img_array[9][14][0] <= img[3744];\
        in_img_array[9][14][1] <= img[3745];\
        in_img_array[9][14][2] <= img[3746];\
        in_img_array[9][14][3] <= img[3747];\
        in_img_array[9][14][4] <= img[3748];\
        in_img_array[9][14][5] <= img[3749];\
        in_img_array[9][14][6] <= img[3750];\
        in_img_array[9][14][7] <= img[3751];\
        in_img_array[9][14][8] <= img[3752];\
        in_img_array[9][14][9] <= img[3753];\
        in_img_array[9][14][10] <= img[3754];\
        in_img_array[9][14][11] <= img[3755];\
        in_img_array[9][14][12] <= img[3756];\
        in_img_array[9][14][13] <= img[3757];\
        in_img_array[9][14][14] <= img[3758];\
        in_img_array[9][14][15] <= img[3759];\
        in_img_array[9][14][16] <= img[3760];\
        in_img_array[9][14][17] <= img[3761];\
        in_img_array[9][15][0] <= img[3762];\
        in_img_array[9][15][1] <= img[3763];\
        in_img_array[9][15][2] <= img[3764];\
        in_img_array[9][15][3] <= img[3765];\
        in_img_array[9][15][4] <= img[3766];\
        in_img_array[9][15][5] <= img[3767];\
        in_img_array[9][15][6] <= img[3768];\
        in_img_array[9][15][7] <= img[3769];\
        in_img_array[9][15][8] <= img[3770];\
        in_img_array[9][15][9] <= img[3771];\
        in_img_array[9][15][10] <= img[3772];\
        in_img_array[9][15][11] <= img[3773];\
        in_img_array[9][15][12] <= img[3774];\
        in_img_array[9][15][13] <= img[3775];\
        in_img_array[9][15][14] <= img[3776];\
        in_img_array[9][15][15] <= img[3777];\
        in_img_array[9][15][16] <= img[3778];\
        in_img_array[9][15][17] <= img[3779];\
        in_img_array[9][16][0] <= img[3780];\
        in_img_array[9][16][1] <= img[3781];\
        in_img_array[9][16][2] <= img[3782];\
        in_img_array[9][16][3] <= img[3783];\
        in_img_array[9][16][4] <= img[3784];\
        in_img_array[9][16][5] <= img[3785];\
        in_img_array[9][16][6] <= img[3786];\
        in_img_array[9][16][7] <= img[3787];\
        in_img_array[9][16][8] <= img[3788];\
        in_img_array[9][16][9] <= img[3789];\
        in_img_array[9][16][10] <= img[3790];\
        in_img_array[9][16][11] <= img[3791];\
        in_img_array[9][16][12] <= img[3792];\
        in_img_array[9][16][13] <= img[3793];\
        in_img_array[9][16][14] <= img[3794];\
        in_img_array[9][16][15] <= img[3795];\
        in_img_array[9][16][16] <= img[3796];\
        in_img_array[9][16][17] <= img[3797];\
        in_img_array[9][17][0] <= img[3798];\
        in_img_array[9][17][1] <= img[3799];\
        in_img_array[9][17][2] <= img[3800];\
        in_img_array[9][17][3] <= img[3801];\
        in_img_array[9][17][4] <= img[3802];\
        in_img_array[9][17][5] <= img[3803];\
        in_img_array[9][17][6] <= img[3804];\
        in_img_array[9][17][7] <= img[3805];\
        in_img_array[9][17][8] <= img[3806];\
        in_img_array[9][17][9] <= img[3807];\
        in_img_array[9][17][10] <= img[3808];\
        in_img_array[9][17][11] <= img[3809];\
        in_img_array[9][17][12] <= img[3810];\
        in_img_array[9][17][13] <= img[3811];\
        in_img_array[9][17][14] <= img[3812];\
        in_img_array[9][17][15] <= img[3813];\
        in_img_array[9][17][16] <= img[3814];\
        in_img_array[9][17][17] <= img[3815];\
        in_img_array[9][18][0] <= img[3816];\
        in_img_array[9][18][1] <= img[3817];\
        in_img_array[9][18][2] <= img[3818];\
        in_img_array[9][18][3] <= img[3819];\
        in_img_array[9][18][4] <= img[3820];\
        in_img_array[9][18][5] <= img[3821];\
        in_img_array[9][18][6] <= img[3822];\
        in_img_array[9][18][7] <= img[3823];\
        in_img_array[9][18][8] <= img[3824];\
        in_img_array[9][18][9] <= img[3825];\
        in_img_array[9][18][10] <= img[3826];\
        in_img_array[9][18][11] <= img[3827];\
        in_img_array[9][18][12] <= img[3828];\
        in_img_array[9][18][13] <= img[3829];\
        in_img_array[9][18][14] <= img[3830];\
        in_img_array[9][18][15] <= img[3831];\
        in_img_array[9][18][16] <= img[3832];\
        in_img_array[9][18][17] <= img[3833];\
        in_img_array[9][19][0] <= img[3834];\
        in_img_array[9][19][1] <= img[3835];\
        in_img_array[9][19][2] <= img[3836];\
        in_img_array[9][19][3] <= img[3837];\
        in_img_array[9][19][4] <= img[3838];\
        in_img_array[9][19][5] <= img[3839];\
        in_img_array[9][19][6] <= img[3840];\
        in_img_array[9][19][7] <= img[3841];\
        in_img_array[9][19][8] <= img[3842];\
        in_img_array[9][19][9] <= img[3843];\
        in_img_array[9][19][10] <= img[3844];\
        in_img_array[9][19][11] <= img[3845];\
        in_img_array[9][19][12] <= img[3846];\
        in_img_array[9][19][13] <= img[3847];\
        in_img_array[9][19][14] <= img[3848];\
        in_img_array[9][19][15] <= img[3849];\
        in_img_array[9][19][16] <= img[3850];\
        in_img_array[9][19][17] <= img[3851];\
        in_img_array[9][20][0] <= img[3852];\
        in_img_array[9][20][1] <= img[3853];\
        in_img_array[9][20][2] <= img[3854];\
        in_img_array[9][20][3] <= img[3855];\
        in_img_array[9][20][4] <= img[3856];\
        in_img_array[9][20][5] <= img[3857];\
        in_img_array[9][20][6] <= img[3858];\
        in_img_array[9][20][7] <= img[3859];\
        in_img_array[9][20][8] <= img[3860];\
        in_img_array[9][20][9] <= img[3861];\
        in_img_array[9][20][10] <= img[3862];\
        in_img_array[9][20][11] <= img[3863];\
        in_img_array[9][20][12] <= img[3864];\
        in_img_array[9][20][13] <= img[3865];\
        in_img_array[9][20][14] <= img[3866];\
        in_img_array[9][20][15] <= img[3867];\
        in_img_array[9][20][16] <= img[3868];\
        in_img_array[9][20][17] <= img[3869];\
        in_img_array[9][21][0] <= img[3870];\
        in_img_array[9][21][1] <= img[3871];\
        in_img_array[9][21][2] <= img[3872];\
        in_img_array[9][21][3] <= img[3873];\
        in_img_array[9][21][4] <= img[3874];\
        in_img_array[9][21][5] <= img[3875];\
        in_img_array[9][21][6] <= img[3876];\
        in_img_array[9][21][7] <= img[3877];\
        in_img_array[9][21][8] <= img[3878];\
        in_img_array[9][21][9] <= img[3879];\
        in_img_array[9][21][10] <= img[3880];\
        in_img_array[9][21][11] <= img[3881];\
        in_img_array[9][21][12] <= img[3882];\
        in_img_array[9][21][13] <= img[3883];\
        in_img_array[9][21][14] <= img[3884];\
        in_img_array[9][21][15] <= img[3885];\
        in_img_array[9][21][16] <= img[3886];\
        in_img_array[9][21][17] <= img[3887];\
        in_img_array[9][22][0] <= img[3888];\
        in_img_array[9][22][1] <= img[3889];\
        in_img_array[9][22][2] <= img[3890];\
        in_img_array[9][22][3] <= img[3891];\
        in_img_array[9][22][4] <= img[3892];\
        in_img_array[9][22][5] <= img[3893];\
        in_img_array[9][22][6] <= img[3894];\
        in_img_array[9][22][7] <= img[3895];\
        in_img_array[9][22][8] <= img[3896];\
        in_img_array[9][22][9] <= img[3897];\
        in_img_array[9][22][10] <= img[3898];\
        in_img_array[9][22][11] <= img[3899];\
        in_img_array[9][22][12] <= img[3900];\
        in_img_array[9][22][13] <= img[3901];\
        in_img_array[9][22][14] <= img[3902];\
        in_img_array[9][22][15] <= img[3903];\
        in_img_array[9][22][16] <= img[3904];\
        in_img_array[9][22][17] <= img[3905];\
        in_img_array[9][23][0] <= img[3906];\
        in_img_array[9][23][1] <= img[3907];\
        in_img_array[9][23][2] <= img[3908];\
        in_img_array[9][23][3] <= img[3909];\
        in_img_array[9][23][4] <= img[3910];\
        in_img_array[9][23][5] <= img[3911];\
        in_img_array[9][23][6] <= img[3912];\
        in_img_array[9][23][7] <= img[3913];\
        in_img_array[9][23][8] <= img[3914];\
        in_img_array[9][23][9] <= img[3915];\
        in_img_array[9][23][10] <= img[3916];\
        in_img_array[9][23][11] <= img[3917];\
        in_img_array[9][23][12] <= img[3918];\
        in_img_array[9][23][13] <= img[3919];\
        in_img_array[9][23][14] <= img[3920];\
        in_img_array[9][23][15] <= img[3921];\
        in_img_array[9][23][16] <= img[3922];\
        in_img_array[9][23][17] <= img[3923];\
        in_img_array[9][24][0] <= img[3924];\
        in_img_array[9][24][1] <= img[3925];\
        in_img_array[9][24][2] <= img[3926];\
        in_img_array[9][24][3] <= img[3927];\
        in_img_array[9][24][4] <= img[3928];\
        in_img_array[9][24][5] <= img[3929];\
        in_img_array[9][24][6] <= img[3930];\
        in_img_array[9][24][7] <= img[3931];\
        in_img_array[9][24][8] <= img[3932];\
        in_img_array[9][24][9] <= img[3933];\
        in_img_array[9][24][10] <= img[3934];\
        in_img_array[9][24][11] <= img[3935];\
        in_img_array[9][24][12] <= img[3936];\
        in_img_array[9][24][13] <= img[3937];\
        in_img_array[9][24][14] <= img[3938];\
        in_img_array[9][24][15] <= img[3939];\
        in_img_array[9][24][16] <= img[3940];\
        in_img_array[9][24][17] <= img[3941];\
        in_img_array[9][25][0] <= img[3942];\
        in_img_array[9][25][1] <= img[3943];\
        in_img_array[9][25][2] <= img[3944];\
        in_img_array[9][25][3] <= img[3945];\
        in_img_array[9][25][4] <= img[3946];\
        in_img_array[9][25][5] <= img[3947];\
        in_img_array[9][25][6] <= img[3948];\
        in_img_array[9][25][7] <= img[3949];\
        in_img_array[9][25][8] <= img[3950];\
        in_img_array[9][25][9] <= img[3951];\
        in_img_array[9][25][10] <= img[3952];\
        in_img_array[9][25][11] <= img[3953];\
        in_img_array[9][25][12] <= img[3954];\
        in_img_array[9][25][13] <= img[3955];\
        in_img_array[9][25][14] <= img[3956];\
        in_img_array[9][25][15] <= img[3957];\
        in_img_array[9][25][16] <= img[3958];\
        in_img_array[9][25][17] <= img[3959];\
        in_img_array[9][26][0] <= img[3960];\
        in_img_array[9][26][1] <= img[3961];\
        in_img_array[9][26][2] <= img[3962];\
        in_img_array[9][26][3] <= img[3963];\
        in_img_array[9][26][4] <= img[3964];\
        in_img_array[9][26][5] <= img[3965];\
        in_img_array[9][26][6] <= img[3966];\
        in_img_array[9][26][7] <= img[3967];\
        in_img_array[9][26][8] <= img[3968];\
        in_img_array[9][26][9] <= img[3969];\
        in_img_array[9][26][10] <= img[3970];\
        in_img_array[9][26][11] <= img[3971];\
        in_img_array[9][26][12] <= img[3972];\
        in_img_array[9][26][13] <= img[3973];\
        in_img_array[9][26][14] <= img[3974];\
        in_img_array[9][26][15] <= img[3975];\
        in_img_array[9][26][16] <= img[3976];\
        in_img_array[9][26][17] <= img[3977];\
        in_img_array[9][27][0] <= img[3978];\
        in_img_array[9][27][1] <= img[3979];\
        in_img_array[9][27][2] <= img[3980];\
        in_img_array[9][27][3] <= img[3981];\
        in_img_array[9][27][4] <= img[3982];\
        in_img_array[9][27][5] <= img[3983];\
        in_img_array[9][27][6] <= img[3984];\
        in_img_array[9][27][7] <= img[3985];\
        in_img_array[9][27][8] <= img[3986];\
        in_img_array[9][27][9] <= img[3987];\
        in_img_array[9][27][10] <= img[3988];\
        in_img_array[9][27][11] <= img[3989];\
        in_img_array[9][27][12] <= img[3990];\
        in_img_array[9][27][13] <= img[3991];\
        in_img_array[9][27][14] <= img[3992];\
        in_img_array[9][27][15] <= img[3993];\
        in_img_array[9][27][16] <= img[3994];\
        in_img_array[9][27][17] <= img[3995];\
        in_img_array[9][28][0] <= img[3996];\
        in_img_array[9][28][1] <= img[3997];\
        in_img_array[9][28][2] <= img[3998];\
        in_img_array[9][28][3] <= img[3999];\
        in_img_array[9][28][4] <= img[4000];\
        in_img_array[9][28][5] <= img[4001];\
        in_img_array[9][28][6] <= img[4002];\
        in_img_array[9][28][7] <= img[4003];\
        in_img_array[9][28][8] <= img[4004];\
        in_img_array[9][28][9] <= img[4005];\
        in_img_array[9][28][10] <= img[4006];\
        in_img_array[9][28][11] <= img[4007];\
        in_img_array[9][28][12] <= img[4008];\
        in_img_array[9][28][13] <= img[4009];\
        in_img_array[9][28][14] <= img[4010];\
        in_img_array[9][28][15] <= img[4011];\
        in_img_array[9][28][16] <= img[4012];\
        in_img_array[9][28][17] <= img[4013];\
        in_img_array[9][29][0] <= img[4014];\
        in_img_array[9][29][1] <= img[4015];\
        in_img_array[9][29][2] <= img[4016];\
        in_img_array[9][29][3] <= img[4017];\
        in_img_array[9][29][4] <= img[4018];\
        in_img_array[9][29][5] <= img[4019];\
        in_img_array[9][29][6] <= img[4020];\
        in_img_array[9][29][7] <= img[4021];\
        in_img_array[9][29][8] <= img[4022];\
        in_img_array[9][29][9] <= img[4023];\
        in_img_array[9][29][10] <= img[4024];\
        in_img_array[9][29][11] <= img[4025];\
        in_img_array[9][29][12] <= img[4026];\
        in_img_array[9][29][13] <= img[4027];\
        in_img_array[9][29][14] <= img[4028];\
        in_img_array[9][29][15] <= img[4029];\
        in_img_array[9][29][16] <= img[4030];\
        in_img_array[9][29][17] <= img[4031];\
        in_img_array[10][2][0] <= img[4032];\
        in_img_array[10][2][1] <= img[4033];\
        in_img_array[10][2][2] <= img[4034];\
        in_img_array[10][2][3] <= img[4035];\
        in_img_array[10][2][4] <= img[4036];\
        in_img_array[10][2][5] <= img[4037];\
        in_img_array[10][2][6] <= img[4038];\
        in_img_array[10][2][7] <= img[4039];\
        in_img_array[10][2][8] <= img[4040];\
        in_img_array[10][2][9] <= img[4041];\
        in_img_array[10][2][10] <= img[4042];\
        in_img_array[10][2][11] <= img[4043];\
        in_img_array[10][2][12] <= img[4044];\
        in_img_array[10][2][13] <= img[4045];\
        in_img_array[10][2][14] <= img[4046];\
        in_img_array[10][2][15] <= img[4047];\
        in_img_array[10][2][16] <= img[4048];\
        in_img_array[10][2][17] <= img[4049];\
        in_img_array[10][3][0] <= img[4050];\
        in_img_array[10][3][1] <= img[4051];\
        in_img_array[10][3][2] <= img[4052];\
        in_img_array[10][3][3] <= img[4053];\
        in_img_array[10][3][4] <= img[4054];\
        in_img_array[10][3][5] <= img[4055];\
        in_img_array[10][3][6] <= img[4056];\
        in_img_array[10][3][7] <= img[4057];\
        in_img_array[10][3][8] <= img[4058];\
        in_img_array[10][3][9] <= img[4059];\
        in_img_array[10][3][10] <= img[4060];\
        in_img_array[10][3][11] <= img[4061];\
        in_img_array[10][3][12] <= img[4062];\
        in_img_array[10][3][13] <= img[4063];\
        in_img_array[10][3][14] <= img[4064];\
        in_img_array[10][3][15] <= img[4065];\
        in_img_array[10][3][16] <= img[4066];\
        in_img_array[10][3][17] <= img[4067];\
        in_img_array[10][4][0] <= img[4068];\
        in_img_array[10][4][1] <= img[4069];\
        in_img_array[10][4][2] <= img[4070];\
        in_img_array[10][4][3] <= img[4071];\
        in_img_array[10][4][4] <= img[4072];\
        in_img_array[10][4][5] <= img[4073];\
        in_img_array[10][4][6] <= img[4074];\
        in_img_array[10][4][7] <= img[4075];\
        in_img_array[10][4][8] <= img[4076];\
        in_img_array[10][4][9] <= img[4077];\
        in_img_array[10][4][10] <= img[4078];\
        in_img_array[10][4][11] <= img[4079];\
        in_img_array[10][4][12] <= img[4080];\
        in_img_array[10][4][13] <= img[4081];\
        in_img_array[10][4][14] <= img[4082];\
        in_img_array[10][4][15] <= img[4083];\
        in_img_array[10][4][16] <= img[4084];\
        in_img_array[10][4][17] <= img[4085];\
        in_img_array[10][5][0] <= img[4086];\
        in_img_array[10][5][1] <= img[4087];\
        in_img_array[10][5][2] <= img[4088];\
        in_img_array[10][5][3] <= img[4089];\
        in_img_array[10][5][4] <= img[4090];\
        in_img_array[10][5][5] <= img[4091];\
        in_img_array[10][5][6] <= img[4092];\
        in_img_array[10][5][7] <= img[4093];\
        in_img_array[10][5][8] <= img[4094];\
        in_img_array[10][5][9] <= img[4095];\
        in_img_array[10][5][10] <= img[4096];\
        in_img_array[10][5][11] <= img[4097];\
        in_img_array[10][5][12] <= img[4098];\
        in_img_array[10][5][13] <= img[4099];\
        in_img_array[10][5][14] <= img[4100];\
        in_img_array[10][5][15] <= img[4101];\
        in_img_array[10][5][16] <= img[4102];\
        in_img_array[10][5][17] <= img[4103];\
        in_img_array[10][6][0] <= img[4104];\
        in_img_array[10][6][1] <= img[4105];\
        in_img_array[10][6][2] <= img[4106];\
        in_img_array[10][6][3] <= img[4107];\
        in_img_array[10][6][4] <= img[4108];\
        in_img_array[10][6][5] <= img[4109];\
        in_img_array[10][6][6] <= img[4110];\
        in_img_array[10][6][7] <= img[4111];\
        in_img_array[10][6][8] <= img[4112];\
        in_img_array[10][6][9] <= img[4113];\
        in_img_array[10][6][10] <= img[4114];\
        in_img_array[10][6][11] <= img[4115];\
        in_img_array[10][6][12] <= img[4116];\
        in_img_array[10][6][13] <= img[4117];\
        in_img_array[10][6][14] <= img[4118];\
        in_img_array[10][6][15] <= img[4119];\
        in_img_array[10][6][16] <= img[4120];\
        in_img_array[10][6][17] <= img[4121];\
        in_img_array[10][7][0] <= img[4122];\
        in_img_array[10][7][1] <= img[4123];\
        in_img_array[10][7][2] <= img[4124];\
        in_img_array[10][7][3] <= img[4125];\
        in_img_array[10][7][4] <= img[4126];\
        in_img_array[10][7][5] <= img[4127];\
        in_img_array[10][7][6] <= img[4128];\
        in_img_array[10][7][7] <= img[4129];\
        in_img_array[10][7][8] <= img[4130];\
        in_img_array[10][7][9] <= img[4131];\
        in_img_array[10][7][10] <= img[4132];\
        in_img_array[10][7][11] <= img[4133];\
        in_img_array[10][7][12] <= img[4134];\
        in_img_array[10][7][13] <= img[4135];\
        in_img_array[10][7][14] <= img[4136];\
        in_img_array[10][7][15] <= img[4137];\
        in_img_array[10][7][16] <= img[4138];\
        in_img_array[10][7][17] <= img[4139];\
        in_img_array[10][8][0] <= img[4140];\
        in_img_array[10][8][1] <= img[4141];\
        in_img_array[10][8][2] <= img[4142];\
        in_img_array[10][8][3] <= img[4143];\
        in_img_array[10][8][4] <= img[4144];\
        in_img_array[10][8][5] <= img[4145];\
        in_img_array[10][8][6] <= img[4146];\
        in_img_array[10][8][7] <= img[4147];\
        in_img_array[10][8][8] <= img[4148];\
        in_img_array[10][8][9] <= img[4149];\
        in_img_array[10][8][10] <= img[4150];\
        in_img_array[10][8][11] <= img[4151];\
        in_img_array[10][8][12] <= img[4152];\
        in_img_array[10][8][13] <= img[4153];\
        in_img_array[10][8][14] <= img[4154];\
        in_img_array[10][8][15] <= img[4155];\
        in_img_array[10][8][16] <= img[4156];\
        in_img_array[10][8][17] <= img[4157];\
        in_img_array[10][9][0] <= img[4158];\
        in_img_array[10][9][1] <= img[4159];\
        in_img_array[10][9][2] <= img[4160];\
        in_img_array[10][9][3] <= img[4161];\
        in_img_array[10][9][4] <= img[4162];\
        in_img_array[10][9][5] <= img[4163];\
        in_img_array[10][9][6] <= img[4164];\
        in_img_array[10][9][7] <= img[4165];\
        in_img_array[10][9][8] <= img[4166];\
        in_img_array[10][9][9] <= img[4167];\
        in_img_array[10][9][10] <= img[4168];\
        in_img_array[10][9][11] <= img[4169];\
        in_img_array[10][9][12] <= img[4170];\
        in_img_array[10][9][13] <= img[4171];\
        in_img_array[10][9][14] <= img[4172];\
        in_img_array[10][9][15] <= img[4173];\
        in_img_array[10][9][16] <= img[4174];\
        in_img_array[10][9][17] <= img[4175];\
        in_img_array[10][10][0] <= img[4176];\
        in_img_array[10][10][1] <= img[4177];\
        in_img_array[10][10][2] <= img[4178];\
        in_img_array[10][10][3] <= img[4179];\
        in_img_array[10][10][4] <= img[4180];\
        in_img_array[10][10][5] <= img[4181];\
        in_img_array[10][10][6] <= img[4182];\
        in_img_array[10][10][7] <= img[4183];\
        in_img_array[10][10][8] <= img[4184];\
        in_img_array[10][10][9] <= img[4185];\
        in_img_array[10][10][10] <= img[4186];\
        in_img_array[10][10][11] <= img[4187];\
        in_img_array[10][10][12] <= img[4188];\
        in_img_array[10][10][13] <= img[4189];\
        in_img_array[10][10][14] <= img[4190];\
        in_img_array[10][10][15] <= img[4191];\
        in_img_array[10][10][16] <= img[4192];\
        in_img_array[10][10][17] <= img[4193];\
        in_img_array[10][11][0] <= img[4194];\
        in_img_array[10][11][1] <= img[4195];\
        in_img_array[10][11][2] <= img[4196];\
        in_img_array[10][11][3] <= img[4197];\
        in_img_array[10][11][4] <= img[4198];\
        in_img_array[10][11][5] <= img[4199];\
        in_img_array[10][11][6] <= img[4200];\
        in_img_array[10][11][7] <= img[4201];\
        in_img_array[10][11][8] <= img[4202];\
        in_img_array[10][11][9] <= img[4203];\
        in_img_array[10][11][10] <= img[4204];\
        in_img_array[10][11][11] <= img[4205];\
        in_img_array[10][11][12] <= img[4206];\
        in_img_array[10][11][13] <= img[4207];\
        in_img_array[10][11][14] <= img[4208];\
        in_img_array[10][11][15] <= img[4209];\
        in_img_array[10][11][16] <= img[4210];\
        in_img_array[10][11][17] <= img[4211];\
        in_img_array[10][12][0] <= img[4212];\
        in_img_array[10][12][1] <= img[4213];\
        in_img_array[10][12][2] <= img[4214];\
        in_img_array[10][12][3] <= img[4215];\
        in_img_array[10][12][4] <= img[4216];\
        in_img_array[10][12][5] <= img[4217];\
        in_img_array[10][12][6] <= img[4218];\
        in_img_array[10][12][7] <= img[4219];\
        in_img_array[10][12][8] <= img[4220];\
        in_img_array[10][12][9] <= img[4221];\
        in_img_array[10][12][10] <= img[4222];\
        in_img_array[10][12][11] <= img[4223];\
        in_img_array[10][12][12] <= img[4224];\
        in_img_array[10][12][13] <= img[4225];\
        in_img_array[10][12][14] <= img[4226];\
        in_img_array[10][12][15] <= img[4227];\
        in_img_array[10][12][16] <= img[4228];\
        in_img_array[10][12][17] <= img[4229];\
        in_img_array[10][13][0] <= img[4230];\
        in_img_array[10][13][1] <= img[4231];\
        in_img_array[10][13][2] <= img[4232];\
        in_img_array[10][13][3] <= img[4233];\
        in_img_array[10][13][4] <= img[4234];\
        in_img_array[10][13][5] <= img[4235];\
        in_img_array[10][13][6] <= img[4236];\
        in_img_array[10][13][7] <= img[4237];\
        in_img_array[10][13][8] <= img[4238];\
        in_img_array[10][13][9] <= img[4239];\
        in_img_array[10][13][10] <= img[4240];\
        in_img_array[10][13][11] <= img[4241];\
        in_img_array[10][13][12] <= img[4242];\
        in_img_array[10][13][13] <= img[4243];\
        in_img_array[10][13][14] <= img[4244];\
        in_img_array[10][13][15] <= img[4245];\
        in_img_array[10][13][16] <= img[4246];\
        in_img_array[10][13][17] <= img[4247];\
        in_img_array[10][14][0] <= img[4248];\
        in_img_array[10][14][1] <= img[4249];\
        in_img_array[10][14][2] <= img[4250];\
        in_img_array[10][14][3] <= img[4251];\
        in_img_array[10][14][4] <= img[4252];\
        in_img_array[10][14][5] <= img[4253];\
        in_img_array[10][14][6] <= img[4254];\
        in_img_array[10][14][7] <= img[4255];\
        in_img_array[10][14][8] <= img[4256];\
        in_img_array[10][14][9] <= img[4257];\
        in_img_array[10][14][10] <= img[4258];\
        in_img_array[10][14][11] <= img[4259];\
        in_img_array[10][14][12] <= img[4260];\
        in_img_array[10][14][13] <= img[4261];\
        in_img_array[10][14][14] <= img[4262];\
        in_img_array[10][14][15] <= img[4263];\
        in_img_array[10][14][16] <= img[4264];\
        in_img_array[10][14][17] <= img[4265];\
        in_img_array[10][15][0] <= img[4266];\
        in_img_array[10][15][1] <= img[4267];\
        in_img_array[10][15][2] <= img[4268];\
        in_img_array[10][15][3] <= img[4269];\
        in_img_array[10][15][4] <= img[4270];\
        in_img_array[10][15][5] <= img[4271];\
        in_img_array[10][15][6] <= img[4272];\
        in_img_array[10][15][7] <= img[4273];\
        in_img_array[10][15][8] <= img[4274];\
        in_img_array[10][15][9] <= img[4275];\
        in_img_array[10][15][10] <= img[4276];\
        in_img_array[10][15][11] <= img[4277];\
        in_img_array[10][15][12] <= img[4278];\
        in_img_array[10][15][13] <= img[4279];\
        in_img_array[10][15][14] <= img[4280];\
        in_img_array[10][15][15] <= img[4281];\
        in_img_array[10][15][16] <= img[4282];\
        in_img_array[10][15][17] <= img[4283];\
        in_img_array[10][16][0] <= img[4284];\
        in_img_array[10][16][1] <= img[4285];\
        in_img_array[10][16][2] <= img[4286];\
        in_img_array[10][16][3] <= img[4287];\
        in_img_array[10][16][4] <= img[4288];\
        in_img_array[10][16][5] <= img[4289];\
        in_img_array[10][16][6] <= img[4290];\
        in_img_array[10][16][7] <= img[4291];\
        in_img_array[10][16][8] <= img[4292];\
        in_img_array[10][16][9] <= img[4293];\
        in_img_array[10][16][10] <= img[4294];\
        in_img_array[10][16][11] <= img[4295];\
        in_img_array[10][16][12] <= img[4296];\
        in_img_array[10][16][13] <= img[4297];\
        in_img_array[10][16][14] <= img[4298];\
        in_img_array[10][16][15] <= img[4299];\
        in_img_array[10][16][16] <= img[4300];\
        in_img_array[10][16][17] <= img[4301];\
        in_img_array[10][17][0] <= img[4302];\
        in_img_array[10][17][1] <= img[4303];\
        in_img_array[10][17][2] <= img[4304];\
        in_img_array[10][17][3] <= img[4305];\
        in_img_array[10][17][4] <= img[4306];\
        in_img_array[10][17][5] <= img[4307];\
        in_img_array[10][17][6] <= img[4308];\
        in_img_array[10][17][7] <= img[4309];\
        in_img_array[10][17][8] <= img[4310];\
        in_img_array[10][17][9] <= img[4311];\
        in_img_array[10][17][10] <= img[4312];\
        in_img_array[10][17][11] <= img[4313];\
        in_img_array[10][17][12] <= img[4314];\
        in_img_array[10][17][13] <= img[4315];\
        in_img_array[10][17][14] <= img[4316];\
        in_img_array[10][17][15] <= img[4317];\
        in_img_array[10][17][16] <= img[4318];\
        in_img_array[10][17][17] <= img[4319];\
        in_img_array[10][18][0] <= img[4320];\
        in_img_array[10][18][1] <= img[4321];\
        in_img_array[10][18][2] <= img[4322];\
        in_img_array[10][18][3] <= img[4323];\
        in_img_array[10][18][4] <= img[4324];\
        in_img_array[10][18][5] <= img[4325];\
        in_img_array[10][18][6] <= img[4326];\
        in_img_array[10][18][7] <= img[4327];\
        in_img_array[10][18][8] <= img[4328];\
        in_img_array[10][18][9] <= img[4329];\
        in_img_array[10][18][10] <= img[4330];\
        in_img_array[10][18][11] <= img[4331];\
        in_img_array[10][18][12] <= img[4332];\
        in_img_array[10][18][13] <= img[4333];\
        in_img_array[10][18][14] <= img[4334];\
        in_img_array[10][18][15] <= img[4335];\
        in_img_array[10][18][16] <= img[4336];\
        in_img_array[10][18][17] <= img[4337];\
        in_img_array[10][19][0] <= img[4338];\
        in_img_array[10][19][1] <= img[4339];\
        in_img_array[10][19][2] <= img[4340];\
        in_img_array[10][19][3] <= img[4341];\
        in_img_array[10][19][4] <= img[4342];\
        in_img_array[10][19][5] <= img[4343];\
        in_img_array[10][19][6] <= img[4344];\
        in_img_array[10][19][7] <= img[4345];\
        in_img_array[10][19][8] <= img[4346];\
        in_img_array[10][19][9] <= img[4347];\
        in_img_array[10][19][10] <= img[4348];\
        in_img_array[10][19][11] <= img[4349];\
        in_img_array[10][19][12] <= img[4350];\
        in_img_array[10][19][13] <= img[4351];\
        in_img_array[10][19][14] <= img[4352];\
        in_img_array[10][19][15] <= img[4353];\
        in_img_array[10][19][16] <= img[4354];\
        in_img_array[10][19][17] <= img[4355];\
        in_img_array[10][20][0] <= img[4356];\
        in_img_array[10][20][1] <= img[4357];\
        in_img_array[10][20][2] <= img[4358];\
        in_img_array[10][20][3] <= img[4359];\
        in_img_array[10][20][4] <= img[4360];\
        in_img_array[10][20][5] <= img[4361];\
        in_img_array[10][20][6] <= img[4362];\
        in_img_array[10][20][7] <= img[4363];\
        in_img_array[10][20][8] <= img[4364];\
        in_img_array[10][20][9] <= img[4365];\
        in_img_array[10][20][10] <= img[4366];\
        in_img_array[10][20][11] <= img[4367];\
        in_img_array[10][20][12] <= img[4368];\
        in_img_array[10][20][13] <= img[4369];\
        in_img_array[10][20][14] <= img[4370];\
        in_img_array[10][20][15] <= img[4371];\
        in_img_array[10][20][16] <= img[4372];\
        in_img_array[10][20][17] <= img[4373];\
        in_img_array[10][21][0] <= img[4374];\
        in_img_array[10][21][1] <= img[4375];\
        in_img_array[10][21][2] <= img[4376];\
        in_img_array[10][21][3] <= img[4377];\
        in_img_array[10][21][4] <= img[4378];\
        in_img_array[10][21][5] <= img[4379];\
        in_img_array[10][21][6] <= img[4380];\
        in_img_array[10][21][7] <= img[4381];\
        in_img_array[10][21][8] <= img[4382];\
        in_img_array[10][21][9] <= img[4383];\
        in_img_array[10][21][10] <= img[4384];\
        in_img_array[10][21][11] <= img[4385];\
        in_img_array[10][21][12] <= img[4386];\
        in_img_array[10][21][13] <= img[4387];\
        in_img_array[10][21][14] <= img[4388];\
        in_img_array[10][21][15] <= img[4389];\
        in_img_array[10][21][16] <= img[4390];\
        in_img_array[10][21][17] <= img[4391];\
        in_img_array[10][22][0] <= img[4392];\
        in_img_array[10][22][1] <= img[4393];\
        in_img_array[10][22][2] <= img[4394];\
        in_img_array[10][22][3] <= img[4395];\
        in_img_array[10][22][4] <= img[4396];\
        in_img_array[10][22][5] <= img[4397];\
        in_img_array[10][22][6] <= img[4398];\
        in_img_array[10][22][7] <= img[4399];\
        in_img_array[10][22][8] <= img[4400];\
        in_img_array[10][22][9] <= img[4401];\
        in_img_array[10][22][10] <= img[4402];\
        in_img_array[10][22][11] <= img[4403];\
        in_img_array[10][22][12] <= img[4404];\
        in_img_array[10][22][13] <= img[4405];\
        in_img_array[10][22][14] <= img[4406];\
        in_img_array[10][22][15] <= img[4407];\
        in_img_array[10][22][16] <= img[4408];\
        in_img_array[10][22][17] <= img[4409];\
        in_img_array[10][23][0] <= img[4410];\
        in_img_array[10][23][1] <= img[4411];\
        in_img_array[10][23][2] <= img[4412];\
        in_img_array[10][23][3] <= img[4413];\
        in_img_array[10][23][4] <= img[4414];\
        in_img_array[10][23][5] <= img[4415];\
        in_img_array[10][23][6] <= img[4416];\
        in_img_array[10][23][7] <= img[4417];\
        in_img_array[10][23][8] <= img[4418];\
        in_img_array[10][23][9] <= img[4419];\
        in_img_array[10][23][10] <= img[4420];\
        in_img_array[10][23][11] <= img[4421];\
        in_img_array[10][23][12] <= img[4422];\
        in_img_array[10][23][13] <= img[4423];\
        in_img_array[10][23][14] <= img[4424];\
        in_img_array[10][23][15] <= img[4425];\
        in_img_array[10][23][16] <= img[4426];\
        in_img_array[10][23][17] <= img[4427];\
        in_img_array[10][24][0] <= img[4428];\
        in_img_array[10][24][1] <= img[4429];\
        in_img_array[10][24][2] <= img[4430];\
        in_img_array[10][24][3] <= img[4431];\
        in_img_array[10][24][4] <= img[4432];\
        in_img_array[10][24][5] <= img[4433];\
        in_img_array[10][24][6] <= img[4434];\
        in_img_array[10][24][7] <= img[4435];\
        in_img_array[10][24][8] <= img[4436];\
        in_img_array[10][24][9] <= img[4437];\
        in_img_array[10][24][10] <= img[4438];\
        in_img_array[10][24][11] <= img[4439];\
        in_img_array[10][24][12] <= img[4440];\
        in_img_array[10][24][13] <= img[4441];\
        in_img_array[10][24][14] <= img[4442];\
        in_img_array[10][24][15] <= img[4443];\
        in_img_array[10][24][16] <= img[4444];\
        in_img_array[10][24][17] <= img[4445];\
        in_img_array[10][25][0] <= img[4446];\
        in_img_array[10][25][1] <= img[4447];\
        in_img_array[10][25][2] <= img[4448];\
        in_img_array[10][25][3] <= img[4449];\
        in_img_array[10][25][4] <= img[4450];\
        in_img_array[10][25][5] <= img[4451];\
        in_img_array[10][25][6] <= img[4452];\
        in_img_array[10][25][7] <= img[4453];\
        in_img_array[10][25][8] <= img[4454];\
        in_img_array[10][25][9] <= img[4455];\
        in_img_array[10][25][10] <= img[4456];\
        in_img_array[10][25][11] <= img[4457];\
        in_img_array[10][25][12] <= img[4458];\
        in_img_array[10][25][13] <= img[4459];\
        in_img_array[10][25][14] <= img[4460];\
        in_img_array[10][25][15] <= img[4461];\
        in_img_array[10][25][16] <= img[4462];\
        in_img_array[10][25][17] <= img[4463];\
        in_img_array[10][26][0] <= img[4464];\
        in_img_array[10][26][1] <= img[4465];\
        in_img_array[10][26][2] <= img[4466];\
        in_img_array[10][26][3] <= img[4467];\
        in_img_array[10][26][4] <= img[4468];\
        in_img_array[10][26][5] <= img[4469];\
        in_img_array[10][26][6] <= img[4470];\
        in_img_array[10][26][7] <= img[4471];\
        in_img_array[10][26][8] <= img[4472];\
        in_img_array[10][26][9] <= img[4473];\
        in_img_array[10][26][10] <= img[4474];\
        in_img_array[10][26][11] <= img[4475];\
        in_img_array[10][26][12] <= img[4476];\
        in_img_array[10][26][13] <= img[4477];\
        in_img_array[10][26][14] <= img[4478];\
        in_img_array[10][26][15] <= img[4479];\
        in_img_array[10][26][16] <= img[4480];\
        in_img_array[10][26][17] <= img[4481];\
        in_img_array[10][27][0] <= img[4482];\
        in_img_array[10][27][1] <= img[4483];\
        in_img_array[10][27][2] <= img[4484];\
        in_img_array[10][27][3] <= img[4485];\
        in_img_array[10][27][4] <= img[4486];\
        in_img_array[10][27][5] <= img[4487];\
        in_img_array[10][27][6] <= img[4488];\
        in_img_array[10][27][7] <= img[4489];\
        in_img_array[10][27][8] <= img[4490];\
        in_img_array[10][27][9] <= img[4491];\
        in_img_array[10][27][10] <= img[4492];\
        in_img_array[10][27][11] <= img[4493];\
        in_img_array[10][27][12] <= img[4494];\
        in_img_array[10][27][13] <= img[4495];\
        in_img_array[10][27][14] <= img[4496];\
        in_img_array[10][27][15] <= img[4497];\
        in_img_array[10][27][16] <= img[4498];\
        in_img_array[10][27][17] <= img[4499];\
        in_img_array[10][28][0] <= img[4500];\
        in_img_array[10][28][1] <= img[4501];\
        in_img_array[10][28][2] <= img[4502];\
        in_img_array[10][28][3] <= img[4503];\
        in_img_array[10][28][4] <= img[4504];\
        in_img_array[10][28][5] <= img[4505];\
        in_img_array[10][28][6] <= img[4506];\
        in_img_array[10][28][7] <= img[4507];\
        in_img_array[10][28][8] <= img[4508];\
        in_img_array[10][28][9] <= img[4509];\
        in_img_array[10][28][10] <= img[4510];\
        in_img_array[10][28][11] <= img[4511];\
        in_img_array[10][28][12] <= img[4512];\
        in_img_array[10][28][13] <= img[4513];\
        in_img_array[10][28][14] <= img[4514];\
        in_img_array[10][28][15] <= img[4515];\
        in_img_array[10][28][16] <= img[4516];\
        in_img_array[10][28][17] <= img[4517];\
        in_img_array[10][29][0] <= img[4518];\
        in_img_array[10][29][1] <= img[4519];\
        in_img_array[10][29][2] <= img[4520];\
        in_img_array[10][29][3] <= img[4521];\
        in_img_array[10][29][4] <= img[4522];\
        in_img_array[10][29][5] <= img[4523];\
        in_img_array[10][29][6] <= img[4524];\
        in_img_array[10][29][7] <= img[4525];\
        in_img_array[10][29][8] <= img[4526];\
        in_img_array[10][29][9] <= img[4527];\
        in_img_array[10][29][10] <= img[4528];\
        in_img_array[10][29][11] <= img[4529];\
        in_img_array[10][29][12] <= img[4530];\
        in_img_array[10][29][13] <= img[4531];\
        in_img_array[10][29][14] <= img[4532];\
        in_img_array[10][29][15] <= img[4533];\
        in_img_array[10][29][16] <= img[4534];\
        in_img_array[10][29][17] <= img[4535];\
        in_img_array[11][2][0] <= img[4536];\
        in_img_array[11][2][1] <= img[4537];\
        in_img_array[11][2][2] <= img[4538];\
        in_img_array[11][2][3] <= img[4539];\
        in_img_array[11][2][4] <= img[4540];\
        in_img_array[11][2][5] <= img[4541];\
        in_img_array[11][2][6] <= img[4542];\
        in_img_array[11][2][7] <= img[4543];\
        in_img_array[11][2][8] <= img[4544];\
        in_img_array[11][2][9] <= img[4545];\
        in_img_array[11][2][10] <= img[4546];\
        in_img_array[11][2][11] <= img[4547];\
        in_img_array[11][2][12] <= img[4548];\
        in_img_array[11][2][13] <= img[4549];\
        in_img_array[11][2][14] <= img[4550];\
        in_img_array[11][2][15] <= img[4551];\
        in_img_array[11][2][16] <= img[4552];\
        in_img_array[11][2][17] <= img[4553];\
        in_img_array[11][3][0] <= img[4554];\
        in_img_array[11][3][1] <= img[4555];\
        in_img_array[11][3][2] <= img[4556];\
        in_img_array[11][3][3] <= img[4557];\
        in_img_array[11][3][4] <= img[4558];\
        in_img_array[11][3][5] <= img[4559];\
        in_img_array[11][3][6] <= img[4560];\
        in_img_array[11][3][7] <= img[4561];\
        in_img_array[11][3][8] <= img[4562];\
        in_img_array[11][3][9] <= img[4563];\
        in_img_array[11][3][10] <= img[4564];\
        in_img_array[11][3][11] <= img[4565];\
        in_img_array[11][3][12] <= img[4566];\
        in_img_array[11][3][13] <= img[4567];\
        in_img_array[11][3][14] <= img[4568];\
        in_img_array[11][3][15] <= img[4569];\
        in_img_array[11][3][16] <= img[4570];\
        in_img_array[11][3][17] <= img[4571];\
        in_img_array[11][4][0] <= img[4572];\
        in_img_array[11][4][1] <= img[4573];\
        in_img_array[11][4][2] <= img[4574];\
        in_img_array[11][4][3] <= img[4575];\
        in_img_array[11][4][4] <= img[4576];\
        in_img_array[11][4][5] <= img[4577];\
        in_img_array[11][4][6] <= img[4578];\
        in_img_array[11][4][7] <= img[4579];\
        in_img_array[11][4][8] <= img[4580];\
        in_img_array[11][4][9] <= img[4581];\
        in_img_array[11][4][10] <= img[4582];\
        in_img_array[11][4][11] <= img[4583];\
        in_img_array[11][4][12] <= img[4584];\
        in_img_array[11][4][13] <= img[4585];\
        in_img_array[11][4][14] <= img[4586];\
        in_img_array[11][4][15] <= img[4587];\
        in_img_array[11][4][16] <= img[4588];\
        in_img_array[11][4][17] <= img[4589];\
        in_img_array[11][5][0] <= img[4590];\
        in_img_array[11][5][1] <= img[4591];\
        in_img_array[11][5][2] <= img[4592];\
        in_img_array[11][5][3] <= img[4593];\
        in_img_array[11][5][4] <= img[4594];\
        in_img_array[11][5][5] <= img[4595];\
        in_img_array[11][5][6] <= img[4596];\
        in_img_array[11][5][7] <= img[4597];\
        in_img_array[11][5][8] <= img[4598];\
        in_img_array[11][5][9] <= img[4599];\
        in_img_array[11][5][10] <= img[4600];\
        in_img_array[11][5][11] <= img[4601];\
        in_img_array[11][5][12] <= img[4602];\
        in_img_array[11][5][13] <= img[4603];\
        in_img_array[11][5][14] <= img[4604];\
        in_img_array[11][5][15] <= img[4605];\
        in_img_array[11][5][16] <= img[4606];\
        in_img_array[11][5][17] <= img[4607];\
        in_img_array[11][6][0] <= img[4608];\
        in_img_array[11][6][1] <= img[4609];\
        in_img_array[11][6][2] <= img[4610];\
        in_img_array[11][6][3] <= img[4611];\
        in_img_array[11][6][4] <= img[4612];\
        in_img_array[11][6][5] <= img[4613];\
        in_img_array[11][6][6] <= img[4614];\
        in_img_array[11][6][7] <= img[4615];\
        in_img_array[11][6][8] <= img[4616];\
        in_img_array[11][6][9] <= img[4617];\
        in_img_array[11][6][10] <= img[4618];\
        in_img_array[11][6][11] <= img[4619];\
        in_img_array[11][6][12] <= img[4620];\
        in_img_array[11][6][13] <= img[4621];\
        in_img_array[11][6][14] <= img[4622];\
        in_img_array[11][6][15] <= img[4623];\
        in_img_array[11][6][16] <= img[4624];\
        in_img_array[11][6][17] <= img[4625];\
        in_img_array[11][7][0] <= img[4626];\
        in_img_array[11][7][1] <= img[4627];\
        in_img_array[11][7][2] <= img[4628];\
        in_img_array[11][7][3] <= img[4629];\
        in_img_array[11][7][4] <= img[4630];\
        in_img_array[11][7][5] <= img[4631];\
        in_img_array[11][7][6] <= img[4632];\
        in_img_array[11][7][7] <= img[4633];\
        in_img_array[11][7][8] <= img[4634];\
        in_img_array[11][7][9] <= img[4635];\
        in_img_array[11][7][10] <= img[4636];\
        in_img_array[11][7][11] <= img[4637];\
        in_img_array[11][7][12] <= img[4638];\
        in_img_array[11][7][13] <= img[4639];\
        in_img_array[11][7][14] <= img[4640];\
        in_img_array[11][7][15] <= img[4641];\
        in_img_array[11][7][16] <= img[4642];\
        in_img_array[11][7][17] <= img[4643];\
        in_img_array[11][8][0] <= img[4644];\
        in_img_array[11][8][1] <= img[4645];\
        in_img_array[11][8][2] <= img[4646];\
        in_img_array[11][8][3] <= img[4647];\
        in_img_array[11][8][4] <= img[4648];\
        in_img_array[11][8][5] <= img[4649];\
        in_img_array[11][8][6] <= img[4650];\
        in_img_array[11][8][7] <= img[4651];\
        in_img_array[11][8][8] <= img[4652];\
        in_img_array[11][8][9] <= img[4653];\
        in_img_array[11][8][10] <= img[4654];\
        in_img_array[11][8][11] <= img[4655];\
        in_img_array[11][8][12] <= img[4656];\
        in_img_array[11][8][13] <= img[4657];\
        in_img_array[11][8][14] <= img[4658];\
        in_img_array[11][8][15] <= img[4659];\
        in_img_array[11][8][16] <= img[4660];\
        in_img_array[11][8][17] <= img[4661];\
        in_img_array[11][9][0] <= img[4662];\
        in_img_array[11][9][1] <= img[4663];\
        in_img_array[11][9][2] <= img[4664];\
        in_img_array[11][9][3] <= img[4665];\
        in_img_array[11][9][4] <= img[4666];\
        in_img_array[11][9][5] <= img[4667];\
        in_img_array[11][9][6] <= img[4668];\
        in_img_array[11][9][7] <= img[4669];\
        in_img_array[11][9][8] <= img[4670];\
        in_img_array[11][9][9] <= img[4671];\
        in_img_array[11][9][10] <= img[4672];\
        in_img_array[11][9][11] <= img[4673];\
        in_img_array[11][9][12] <= img[4674];\
        in_img_array[11][9][13] <= img[4675];\
        in_img_array[11][9][14] <= img[4676];\
        in_img_array[11][9][15] <= img[4677];\
        in_img_array[11][9][16] <= img[4678];\
        in_img_array[11][9][17] <= img[4679];\
        in_img_array[11][10][0] <= img[4680];\
        in_img_array[11][10][1] <= img[4681];\
        in_img_array[11][10][2] <= img[4682];\
        in_img_array[11][10][3] <= img[4683];\
        in_img_array[11][10][4] <= img[4684];\
        in_img_array[11][10][5] <= img[4685];\
        in_img_array[11][10][6] <= img[4686];\
        in_img_array[11][10][7] <= img[4687];\
        in_img_array[11][10][8] <= img[4688];\
        in_img_array[11][10][9] <= img[4689];\
        in_img_array[11][10][10] <= img[4690];\
        in_img_array[11][10][11] <= img[4691];\
        in_img_array[11][10][12] <= img[4692];\
        in_img_array[11][10][13] <= img[4693];\
        in_img_array[11][10][14] <= img[4694];\
        in_img_array[11][10][15] <= img[4695];\
        in_img_array[11][10][16] <= img[4696];\
        in_img_array[11][10][17] <= img[4697];\
        in_img_array[11][11][0] <= img[4698];\
        in_img_array[11][11][1] <= img[4699];\
        in_img_array[11][11][2] <= img[4700];\
        in_img_array[11][11][3] <= img[4701];\
        in_img_array[11][11][4] <= img[4702];\
        in_img_array[11][11][5] <= img[4703];\
        in_img_array[11][11][6] <= img[4704];\
        in_img_array[11][11][7] <= img[4705];\
        in_img_array[11][11][8] <= img[4706];\
        in_img_array[11][11][9] <= img[4707];\
        in_img_array[11][11][10] <= img[4708];\
        in_img_array[11][11][11] <= img[4709];\
        in_img_array[11][11][12] <= img[4710];\
        in_img_array[11][11][13] <= img[4711];\
        in_img_array[11][11][14] <= img[4712];\
        in_img_array[11][11][15] <= img[4713];\
        in_img_array[11][11][16] <= img[4714];\
        in_img_array[11][11][17] <= img[4715];\
        in_img_array[11][12][0] <= img[4716];\
        in_img_array[11][12][1] <= img[4717];\
        in_img_array[11][12][2] <= img[4718];\
        in_img_array[11][12][3] <= img[4719];\
        in_img_array[11][12][4] <= img[4720];\
        in_img_array[11][12][5] <= img[4721];\
        in_img_array[11][12][6] <= img[4722];\
        in_img_array[11][12][7] <= img[4723];\
        in_img_array[11][12][8] <= img[4724];\
        in_img_array[11][12][9] <= img[4725];\
        in_img_array[11][12][10] <= img[4726];\
        in_img_array[11][12][11] <= img[4727];\
        in_img_array[11][12][12] <= img[4728];\
        in_img_array[11][12][13] <= img[4729];\
        in_img_array[11][12][14] <= img[4730];\
        in_img_array[11][12][15] <= img[4731];\
        in_img_array[11][12][16] <= img[4732];\
        in_img_array[11][12][17] <= img[4733];\
        in_img_array[11][13][0] <= img[4734];\
        in_img_array[11][13][1] <= img[4735];\
        in_img_array[11][13][2] <= img[4736];\
        in_img_array[11][13][3] <= img[4737];\
        in_img_array[11][13][4] <= img[4738];\
        in_img_array[11][13][5] <= img[4739];\
        in_img_array[11][13][6] <= img[4740];\
        in_img_array[11][13][7] <= img[4741];\
        in_img_array[11][13][8] <= img[4742];\
        in_img_array[11][13][9] <= img[4743];\
        in_img_array[11][13][10] <= img[4744];\
        in_img_array[11][13][11] <= img[4745];\
        in_img_array[11][13][12] <= img[4746];\
        in_img_array[11][13][13] <= img[4747];\
        in_img_array[11][13][14] <= img[4748];\
        in_img_array[11][13][15] <= img[4749];\
        in_img_array[11][13][16] <= img[4750];\
        in_img_array[11][13][17] <= img[4751];\
        in_img_array[11][14][0] <= img[4752];\
        in_img_array[11][14][1] <= img[4753];\
        in_img_array[11][14][2] <= img[4754];\
        in_img_array[11][14][3] <= img[4755];\
        in_img_array[11][14][4] <= img[4756];\
        in_img_array[11][14][5] <= img[4757];\
        in_img_array[11][14][6] <= img[4758];\
        in_img_array[11][14][7] <= img[4759];\
        in_img_array[11][14][8] <= img[4760];\
        in_img_array[11][14][9] <= img[4761];\
        in_img_array[11][14][10] <= img[4762];\
        in_img_array[11][14][11] <= img[4763];\
        in_img_array[11][14][12] <= img[4764];\
        in_img_array[11][14][13] <= img[4765];\
        in_img_array[11][14][14] <= img[4766];\
        in_img_array[11][14][15] <= img[4767];\
        in_img_array[11][14][16] <= img[4768];\
        in_img_array[11][14][17] <= img[4769];\
        in_img_array[11][15][0] <= img[4770];\
        in_img_array[11][15][1] <= img[4771];\
        in_img_array[11][15][2] <= img[4772];\
        in_img_array[11][15][3] <= img[4773];\
        in_img_array[11][15][4] <= img[4774];\
        in_img_array[11][15][5] <= img[4775];\
        in_img_array[11][15][6] <= img[4776];\
        in_img_array[11][15][7] <= img[4777];\
        in_img_array[11][15][8] <= img[4778];\
        in_img_array[11][15][9] <= img[4779];\
        in_img_array[11][15][10] <= img[4780];\
        in_img_array[11][15][11] <= img[4781];\
        in_img_array[11][15][12] <= img[4782];\
        in_img_array[11][15][13] <= img[4783];\
        in_img_array[11][15][14] <= img[4784];\
        in_img_array[11][15][15] <= img[4785];\
        in_img_array[11][15][16] <= img[4786];\
        in_img_array[11][15][17] <= img[4787];\
        in_img_array[11][16][0] <= img[4788];\
        in_img_array[11][16][1] <= img[4789];\
        in_img_array[11][16][2] <= img[4790];\
        in_img_array[11][16][3] <= img[4791];\
        in_img_array[11][16][4] <= img[4792];\
        in_img_array[11][16][5] <= img[4793];\
        in_img_array[11][16][6] <= img[4794];\
        in_img_array[11][16][7] <= img[4795];\
        in_img_array[11][16][8] <= img[4796];\
        in_img_array[11][16][9] <= img[4797];\
        in_img_array[11][16][10] <= img[4798];\
        in_img_array[11][16][11] <= img[4799];\
        in_img_array[11][16][12] <= img[4800];\
        in_img_array[11][16][13] <= img[4801];\
        in_img_array[11][16][14] <= img[4802];\
        in_img_array[11][16][15] <= img[4803];\
        in_img_array[11][16][16] <= img[4804];\
        in_img_array[11][16][17] <= img[4805];\
        in_img_array[11][17][0] <= img[4806];\
        in_img_array[11][17][1] <= img[4807];\
        in_img_array[11][17][2] <= img[4808];\
        in_img_array[11][17][3] <= img[4809];\
        in_img_array[11][17][4] <= img[4810];\
        in_img_array[11][17][5] <= img[4811];\
        in_img_array[11][17][6] <= img[4812];\
        in_img_array[11][17][7] <= img[4813];\
        in_img_array[11][17][8] <= img[4814];\
        in_img_array[11][17][9] <= img[4815];\
        in_img_array[11][17][10] <= img[4816];\
        in_img_array[11][17][11] <= img[4817];\
        in_img_array[11][17][12] <= img[4818];\
        in_img_array[11][17][13] <= img[4819];\
        in_img_array[11][17][14] <= img[4820];\
        in_img_array[11][17][15] <= img[4821];\
        in_img_array[11][17][16] <= img[4822];\
        in_img_array[11][17][17] <= img[4823];\
        in_img_array[11][18][0] <= img[4824];\
        in_img_array[11][18][1] <= img[4825];\
        in_img_array[11][18][2] <= img[4826];\
        in_img_array[11][18][3] <= img[4827];\
        in_img_array[11][18][4] <= img[4828];\
        in_img_array[11][18][5] <= img[4829];\
        in_img_array[11][18][6] <= img[4830];\
        in_img_array[11][18][7] <= img[4831];\
        in_img_array[11][18][8] <= img[4832];\
        in_img_array[11][18][9] <= img[4833];\
        in_img_array[11][18][10] <= img[4834];\
        in_img_array[11][18][11] <= img[4835];\
        in_img_array[11][18][12] <= img[4836];\
        in_img_array[11][18][13] <= img[4837];\
        in_img_array[11][18][14] <= img[4838];\
        in_img_array[11][18][15] <= img[4839];\
        in_img_array[11][18][16] <= img[4840];\
        in_img_array[11][18][17] <= img[4841];\
        in_img_array[11][19][0] <= img[4842];\
        in_img_array[11][19][1] <= img[4843];\
        in_img_array[11][19][2] <= img[4844];\
        in_img_array[11][19][3] <= img[4845];\
        in_img_array[11][19][4] <= img[4846];\
        in_img_array[11][19][5] <= img[4847];\
        in_img_array[11][19][6] <= img[4848];\
        in_img_array[11][19][7] <= img[4849];\
        in_img_array[11][19][8] <= img[4850];\
        in_img_array[11][19][9] <= img[4851];\
        in_img_array[11][19][10] <= img[4852];\
        in_img_array[11][19][11] <= img[4853];\
        in_img_array[11][19][12] <= img[4854];\
        in_img_array[11][19][13] <= img[4855];\
        in_img_array[11][19][14] <= img[4856];\
        in_img_array[11][19][15] <= img[4857];\
        in_img_array[11][19][16] <= img[4858];\
        in_img_array[11][19][17] <= img[4859];\
        in_img_array[11][20][0] <= img[4860];\
        in_img_array[11][20][1] <= img[4861];\
        in_img_array[11][20][2] <= img[4862];\
        in_img_array[11][20][3] <= img[4863];\
        in_img_array[11][20][4] <= img[4864];\
        in_img_array[11][20][5] <= img[4865];\
        in_img_array[11][20][6] <= img[4866];\
        in_img_array[11][20][7] <= img[4867];\
        in_img_array[11][20][8] <= img[4868];\
        in_img_array[11][20][9] <= img[4869];\
        in_img_array[11][20][10] <= img[4870];\
        in_img_array[11][20][11] <= img[4871];\
        in_img_array[11][20][12] <= img[4872];\
        in_img_array[11][20][13] <= img[4873];\
        in_img_array[11][20][14] <= img[4874];\
        in_img_array[11][20][15] <= img[4875];\
        in_img_array[11][20][16] <= img[4876];\
        in_img_array[11][20][17] <= img[4877];\
        in_img_array[11][21][0] <= img[4878];\
        in_img_array[11][21][1] <= img[4879];\
        in_img_array[11][21][2] <= img[4880];\
        in_img_array[11][21][3] <= img[4881];\
        in_img_array[11][21][4] <= img[4882];\
        in_img_array[11][21][5] <= img[4883];\
        in_img_array[11][21][6] <= img[4884];\
        in_img_array[11][21][7] <= img[4885];\
        in_img_array[11][21][8] <= img[4886];\
        in_img_array[11][21][9] <= img[4887];\
        in_img_array[11][21][10] <= img[4888];\
        in_img_array[11][21][11] <= img[4889];\
        in_img_array[11][21][12] <= img[4890];\
        in_img_array[11][21][13] <= img[4891];\
        in_img_array[11][21][14] <= img[4892];\
        in_img_array[11][21][15] <= img[4893];\
        in_img_array[11][21][16] <= img[4894];\
        in_img_array[11][21][17] <= img[4895];\
        in_img_array[11][22][0] <= img[4896];\
        in_img_array[11][22][1] <= img[4897];\
        in_img_array[11][22][2] <= img[4898];\
        in_img_array[11][22][3] <= img[4899];\
        in_img_array[11][22][4] <= img[4900];\
        in_img_array[11][22][5] <= img[4901];\
        in_img_array[11][22][6] <= img[4902];\
        in_img_array[11][22][7] <= img[4903];\
        in_img_array[11][22][8] <= img[4904];\
        in_img_array[11][22][9] <= img[4905];\
        in_img_array[11][22][10] <= img[4906];\
        in_img_array[11][22][11] <= img[4907];\
        in_img_array[11][22][12] <= img[4908];\
        in_img_array[11][22][13] <= img[4909];\
        in_img_array[11][22][14] <= img[4910];\
        in_img_array[11][22][15] <= img[4911];\
        in_img_array[11][22][16] <= img[4912];\
        in_img_array[11][22][17] <= img[4913];\
        in_img_array[11][23][0] <= img[4914];\
        in_img_array[11][23][1] <= img[4915];\
        in_img_array[11][23][2] <= img[4916];\
        in_img_array[11][23][3] <= img[4917];\
        in_img_array[11][23][4] <= img[4918];\
        in_img_array[11][23][5] <= img[4919];\
        in_img_array[11][23][6] <= img[4920];\
        in_img_array[11][23][7] <= img[4921];\
        in_img_array[11][23][8] <= img[4922];\
        in_img_array[11][23][9] <= img[4923];\
        in_img_array[11][23][10] <= img[4924];\
        in_img_array[11][23][11] <= img[4925];\
        in_img_array[11][23][12] <= img[4926];\
        in_img_array[11][23][13] <= img[4927];\
        in_img_array[11][23][14] <= img[4928];\
        in_img_array[11][23][15] <= img[4929];\
        in_img_array[11][23][16] <= img[4930];\
        in_img_array[11][23][17] <= img[4931];\
        in_img_array[11][24][0] <= img[4932];\
        in_img_array[11][24][1] <= img[4933];\
        in_img_array[11][24][2] <= img[4934];\
        in_img_array[11][24][3] <= img[4935];\
        in_img_array[11][24][4] <= img[4936];\
        in_img_array[11][24][5] <= img[4937];\
        in_img_array[11][24][6] <= img[4938];\
        in_img_array[11][24][7] <= img[4939];\
        in_img_array[11][24][8] <= img[4940];\
        in_img_array[11][24][9] <= img[4941];\
        in_img_array[11][24][10] <= img[4942];\
        in_img_array[11][24][11] <= img[4943];\
        in_img_array[11][24][12] <= img[4944];\
        in_img_array[11][24][13] <= img[4945];\
        in_img_array[11][24][14] <= img[4946];\
        in_img_array[11][24][15] <= img[4947];\
        in_img_array[11][24][16] <= img[4948];\
        in_img_array[11][24][17] <= img[4949];\
        in_img_array[11][25][0] <= img[4950];\
        in_img_array[11][25][1] <= img[4951];\
        in_img_array[11][25][2] <= img[4952];\
        in_img_array[11][25][3] <= img[4953];\
        in_img_array[11][25][4] <= img[4954];\
        in_img_array[11][25][5] <= img[4955];\
        in_img_array[11][25][6] <= img[4956];\
        in_img_array[11][25][7] <= img[4957];\
        in_img_array[11][25][8] <= img[4958];\
        in_img_array[11][25][9] <= img[4959];\
        in_img_array[11][25][10] <= img[4960];\
        in_img_array[11][25][11] <= img[4961];\
        in_img_array[11][25][12] <= img[4962];\
        in_img_array[11][25][13] <= img[4963];\
        in_img_array[11][25][14] <= img[4964];\
        in_img_array[11][25][15] <= img[4965];\
        in_img_array[11][25][16] <= img[4966];\
        in_img_array[11][25][17] <= img[4967];\
        in_img_array[11][26][0] <= img[4968];\
        in_img_array[11][26][1] <= img[4969];\
        in_img_array[11][26][2] <= img[4970];\
        in_img_array[11][26][3] <= img[4971];\
        in_img_array[11][26][4] <= img[4972];\
        in_img_array[11][26][5] <= img[4973];\
        in_img_array[11][26][6] <= img[4974];\
        in_img_array[11][26][7] <= img[4975];\
        in_img_array[11][26][8] <= img[4976];\
        in_img_array[11][26][9] <= img[4977];\
        in_img_array[11][26][10] <= img[4978];\
        in_img_array[11][26][11] <= img[4979];\
        in_img_array[11][26][12] <= img[4980];\
        in_img_array[11][26][13] <= img[4981];\
        in_img_array[11][26][14] <= img[4982];\
        in_img_array[11][26][15] <= img[4983];\
        in_img_array[11][26][16] <= img[4984];\
        in_img_array[11][26][17] <= img[4985];\
        in_img_array[11][27][0] <= img[4986];\
        in_img_array[11][27][1] <= img[4987];\
        in_img_array[11][27][2] <= img[4988];\
        in_img_array[11][27][3] <= img[4989];\
        in_img_array[11][27][4] <= img[4990];\
        in_img_array[11][27][5] <= img[4991];\
        in_img_array[11][27][6] <= img[4992];\
        in_img_array[11][27][7] <= img[4993];\
        in_img_array[11][27][8] <= img[4994];\
        in_img_array[11][27][9] <= img[4995];\
        in_img_array[11][27][10] <= img[4996];\
        in_img_array[11][27][11] <= img[4997];\
        in_img_array[11][27][12] <= img[4998];\
        in_img_array[11][27][13] <= img[4999];\
        in_img_array[11][27][14] <= img[5000];\
        in_img_array[11][27][15] <= img[5001];\
        in_img_array[11][27][16] <= img[5002];\
        in_img_array[11][27][17] <= img[5003];\
        in_img_array[11][28][0] <= img[5004];\
        in_img_array[11][28][1] <= img[5005];\
        in_img_array[11][28][2] <= img[5006];\
        in_img_array[11][28][3] <= img[5007];\
        in_img_array[11][28][4] <= img[5008];\
        in_img_array[11][28][5] <= img[5009];\
        in_img_array[11][28][6] <= img[5010];\
        in_img_array[11][28][7] <= img[5011];\
        in_img_array[11][28][8] <= img[5012];\
        in_img_array[11][28][9] <= img[5013];\
        in_img_array[11][28][10] <= img[5014];\
        in_img_array[11][28][11] <= img[5015];\
        in_img_array[11][28][12] <= img[5016];\
        in_img_array[11][28][13] <= img[5017];\
        in_img_array[11][28][14] <= img[5018];\
        in_img_array[11][28][15] <= img[5019];\
        in_img_array[11][28][16] <= img[5020];\
        in_img_array[11][28][17] <= img[5021];\
        in_img_array[11][29][0] <= img[5022];\
        in_img_array[11][29][1] <= img[5023];\
        in_img_array[11][29][2] <= img[5024];\
        in_img_array[11][29][3] <= img[5025];\
        in_img_array[11][29][4] <= img[5026];\
        in_img_array[11][29][5] <= img[5027];\
        in_img_array[11][29][6] <= img[5028];\
        in_img_array[11][29][7] <= img[5029];\
        in_img_array[11][29][8] <= img[5030];\
        in_img_array[11][29][9] <= img[5031];\
        in_img_array[11][29][10] <= img[5032];\
        in_img_array[11][29][11] <= img[5033];\
        in_img_array[11][29][12] <= img[5034];\
        in_img_array[11][29][13] <= img[5035];\
        in_img_array[11][29][14] <= img[5036];\
        in_img_array[11][29][15] <= img[5037];\
        in_img_array[11][29][16] <= img[5038];\
        in_img_array[11][29][17] <= img[5039];\
        in_img_array[12][2][0] <= img[5040];\
        in_img_array[12][2][1] <= img[5041];\
        in_img_array[12][2][2] <= img[5042];\
        in_img_array[12][2][3] <= img[5043];\
        in_img_array[12][2][4] <= img[5044];\
        in_img_array[12][2][5] <= img[5045];\
        in_img_array[12][2][6] <= img[5046];\
        in_img_array[12][2][7] <= img[5047];\
        in_img_array[12][2][8] <= img[5048];\
        in_img_array[12][2][9] <= img[5049];\
        in_img_array[12][2][10] <= img[5050];\
        in_img_array[12][2][11] <= img[5051];\
        in_img_array[12][2][12] <= img[5052];\
        in_img_array[12][2][13] <= img[5053];\
        in_img_array[12][2][14] <= img[5054];\
        in_img_array[12][2][15] <= img[5055];\
        in_img_array[12][2][16] <= img[5056];\
        in_img_array[12][2][17] <= img[5057];\
        in_img_array[12][3][0] <= img[5058];\
        in_img_array[12][3][1] <= img[5059];\
        in_img_array[12][3][2] <= img[5060];\
        in_img_array[12][3][3] <= img[5061];\
        in_img_array[12][3][4] <= img[5062];\
        in_img_array[12][3][5] <= img[5063];\
        in_img_array[12][3][6] <= img[5064];\
        in_img_array[12][3][7] <= img[5065];\
        in_img_array[12][3][8] <= img[5066];\
        in_img_array[12][3][9] <= img[5067];\
        in_img_array[12][3][10] <= img[5068];\
        in_img_array[12][3][11] <= img[5069];\
        in_img_array[12][3][12] <= img[5070];\
        in_img_array[12][3][13] <= img[5071];\
        in_img_array[12][3][14] <= img[5072];\
        in_img_array[12][3][15] <= img[5073];\
        in_img_array[12][3][16] <= img[5074];\
        in_img_array[12][3][17] <= img[5075];\
        in_img_array[12][4][0] <= img[5076];\
        in_img_array[12][4][1] <= img[5077];\
        in_img_array[12][4][2] <= img[5078];\
        in_img_array[12][4][3] <= img[5079];\
        in_img_array[12][4][4] <= img[5080];\
        in_img_array[12][4][5] <= img[5081];\
        in_img_array[12][4][6] <= img[5082];\
        in_img_array[12][4][7] <= img[5083];\
        in_img_array[12][4][8] <= img[5084];\
        in_img_array[12][4][9] <= img[5085];\
        in_img_array[12][4][10] <= img[5086];\
        in_img_array[12][4][11] <= img[5087];\
        in_img_array[12][4][12] <= img[5088];\
        in_img_array[12][4][13] <= img[5089];\
        in_img_array[12][4][14] <= img[5090];\
        in_img_array[12][4][15] <= img[5091];\
        in_img_array[12][4][16] <= img[5092];\
        in_img_array[12][4][17] <= img[5093];\
        in_img_array[12][5][0] <= img[5094];\
        in_img_array[12][5][1] <= img[5095];\
        in_img_array[12][5][2] <= img[5096];\
        in_img_array[12][5][3] <= img[5097];\
        in_img_array[12][5][4] <= img[5098];\
        in_img_array[12][5][5] <= img[5099];\
        in_img_array[12][5][6] <= img[5100];\
        in_img_array[12][5][7] <= img[5101];\
        in_img_array[12][5][8] <= img[5102];\
        in_img_array[12][5][9] <= img[5103];\
        in_img_array[12][5][10] <= img[5104];\
        in_img_array[12][5][11] <= img[5105];\
        in_img_array[12][5][12] <= img[5106];\
        in_img_array[12][5][13] <= img[5107];\
        in_img_array[12][5][14] <= img[5108];\
        in_img_array[12][5][15] <= img[5109];\
        in_img_array[12][5][16] <= img[5110];\
        in_img_array[12][5][17] <= img[5111];\
        in_img_array[12][6][0] <= img[5112];\
        in_img_array[12][6][1] <= img[5113];\
        in_img_array[12][6][2] <= img[5114];\
        in_img_array[12][6][3] <= img[5115];\
        in_img_array[12][6][4] <= img[5116];\
        in_img_array[12][6][5] <= img[5117];\
        in_img_array[12][6][6] <= img[5118];\
        in_img_array[12][6][7] <= img[5119];\
        in_img_array[12][6][8] <= img[5120];\
        in_img_array[12][6][9] <= img[5121];\
        in_img_array[12][6][10] <= img[5122];\
        in_img_array[12][6][11] <= img[5123];\
        in_img_array[12][6][12] <= img[5124];\
        in_img_array[12][6][13] <= img[5125];\
        in_img_array[12][6][14] <= img[5126];\
        in_img_array[12][6][15] <= img[5127];\
        in_img_array[12][6][16] <= img[5128];\
        in_img_array[12][6][17] <= img[5129];\
        in_img_array[12][7][0] <= img[5130];\
        in_img_array[12][7][1] <= img[5131];\
        in_img_array[12][7][2] <= img[5132];\
        in_img_array[12][7][3] <= img[5133];\
        in_img_array[12][7][4] <= img[5134];\
        in_img_array[12][7][5] <= img[5135];\
        in_img_array[12][7][6] <= img[5136];\
        in_img_array[12][7][7] <= img[5137];\
        in_img_array[12][7][8] <= img[5138];\
        in_img_array[12][7][9] <= img[5139];\
        in_img_array[12][7][10] <= img[5140];\
        in_img_array[12][7][11] <= img[5141];\
        in_img_array[12][7][12] <= img[5142];\
        in_img_array[12][7][13] <= img[5143];\
        in_img_array[12][7][14] <= img[5144];\
        in_img_array[12][7][15] <= img[5145];\
        in_img_array[12][7][16] <= img[5146];\
        in_img_array[12][7][17] <= img[5147];\
        in_img_array[12][8][0] <= img[5148];\
        in_img_array[12][8][1] <= img[5149];\
        in_img_array[12][8][2] <= img[5150];\
        in_img_array[12][8][3] <= img[5151];\
        in_img_array[12][8][4] <= img[5152];\
        in_img_array[12][8][5] <= img[5153];\
        in_img_array[12][8][6] <= img[5154];\
        in_img_array[12][8][7] <= img[5155];\
        in_img_array[12][8][8] <= img[5156];\
        in_img_array[12][8][9] <= img[5157];\
        in_img_array[12][8][10] <= img[5158];\
        in_img_array[12][8][11] <= img[5159];\
        in_img_array[12][8][12] <= img[5160];\
        in_img_array[12][8][13] <= img[5161];\
        in_img_array[12][8][14] <= img[5162];\
        in_img_array[12][8][15] <= img[5163];\
        in_img_array[12][8][16] <= img[5164];\
        in_img_array[12][8][17] <= img[5165];\
        in_img_array[12][9][0] <= img[5166];\
        in_img_array[12][9][1] <= img[5167];\
        in_img_array[12][9][2] <= img[5168];\
        in_img_array[12][9][3] <= img[5169];\
        in_img_array[12][9][4] <= img[5170];\
        in_img_array[12][9][5] <= img[5171];\
        in_img_array[12][9][6] <= img[5172];\
        in_img_array[12][9][7] <= img[5173];\
        in_img_array[12][9][8] <= img[5174];\
        in_img_array[12][9][9] <= img[5175];\
        in_img_array[12][9][10] <= img[5176];\
        in_img_array[12][9][11] <= img[5177];\
        in_img_array[12][9][12] <= img[5178];\
        in_img_array[12][9][13] <= img[5179];\
        in_img_array[12][9][14] <= img[5180];\
        in_img_array[12][9][15] <= img[5181];\
        in_img_array[12][9][16] <= img[5182];\
        in_img_array[12][9][17] <= img[5183];\
        in_img_array[12][10][0] <= img[5184];\
        in_img_array[12][10][1] <= img[5185];\
        in_img_array[12][10][2] <= img[5186];\
        in_img_array[12][10][3] <= img[5187];\
        in_img_array[12][10][4] <= img[5188];\
        in_img_array[12][10][5] <= img[5189];\
        in_img_array[12][10][6] <= img[5190];\
        in_img_array[12][10][7] <= img[5191];\
        in_img_array[12][10][8] <= img[5192];\
        in_img_array[12][10][9] <= img[5193];\
        in_img_array[12][10][10] <= img[5194];\
        in_img_array[12][10][11] <= img[5195];\
        in_img_array[12][10][12] <= img[5196];\
        in_img_array[12][10][13] <= img[5197];\
        in_img_array[12][10][14] <= img[5198];\
        in_img_array[12][10][15] <= img[5199];\
        in_img_array[12][10][16] <= img[5200];\
        in_img_array[12][10][17] <= img[5201];\
        in_img_array[12][11][0] <= img[5202];\
        in_img_array[12][11][1] <= img[5203];\
        in_img_array[12][11][2] <= img[5204];\
        in_img_array[12][11][3] <= img[5205];\
        in_img_array[12][11][4] <= img[5206];\
        in_img_array[12][11][5] <= img[5207];\
        in_img_array[12][11][6] <= img[5208];\
        in_img_array[12][11][7] <= img[5209];\
        in_img_array[12][11][8] <= img[5210];\
        in_img_array[12][11][9] <= img[5211];\
        in_img_array[12][11][10] <= img[5212];\
        in_img_array[12][11][11] <= img[5213];\
        in_img_array[12][11][12] <= img[5214];\
        in_img_array[12][11][13] <= img[5215];\
        in_img_array[12][11][14] <= img[5216];\
        in_img_array[12][11][15] <= img[5217];\
        in_img_array[12][11][16] <= img[5218];\
        in_img_array[12][11][17] <= img[5219];\
        in_img_array[12][12][0] <= img[5220];\
        in_img_array[12][12][1] <= img[5221];\
        in_img_array[12][12][2] <= img[5222];\
        in_img_array[12][12][3] <= img[5223];\
        in_img_array[12][12][4] <= img[5224];\
        in_img_array[12][12][5] <= img[5225];\
        in_img_array[12][12][6] <= img[5226];\
        in_img_array[12][12][7] <= img[5227];\
        in_img_array[12][12][8] <= img[5228];\
        in_img_array[12][12][9] <= img[5229];\
        in_img_array[12][12][10] <= img[5230];\
        in_img_array[12][12][11] <= img[5231];\
        in_img_array[12][12][12] <= img[5232];\
        in_img_array[12][12][13] <= img[5233];\
        in_img_array[12][12][14] <= img[5234];\
        in_img_array[12][12][15] <= img[5235];\
        in_img_array[12][12][16] <= img[5236];\
        in_img_array[12][12][17] <= img[5237];\
        in_img_array[12][13][0] <= img[5238];\
        in_img_array[12][13][1] <= img[5239];\
        in_img_array[12][13][2] <= img[5240];\
        in_img_array[12][13][3] <= img[5241];\
        in_img_array[12][13][4] <= img[5242];\
        in_img_array[12][13][5] <= img[5243];\
        in_img_array[12][13][6] <= img[5244];\
        in_img_array[12][13][7] <= img[5245];\
        in_img_array[12][13][8] <= img[5246];\
        in_img_array[12][13][9] <= img[5247];\
        in_img_array[12][13][10] <= img[5248];\
        in_img_array[12][13][11] <= img[5249];\
        in_img_array[12][13][12] <= img[5250];\
        in_img_array[12][13][13] <= img[5251];\
        in_img_array[12][13][14] <= img[5252];\
        in_img_array[12][13][15] <= img[5253];\
        in_img_array[12][13][16] <= img[5254];\
        in_img_array[12][13][17] <= img[5255];\
        in_img_array[12][14][0] <= img[5256];\
        in_img_array[12][14][1] <= img[5257];\
        in_img_array[12][14][2] <= img[5258];\
        in_img_array[12][14][3] <= img[5259];\
        in_img_array[12][14][4] <= img[5260];\
        in_img_array[12][14][5] <= img[5261];\
        in_img_array[12][14][6] <= img[5262];\
        in_img_array[12][14][7] <= img[5263];\
        in_img_array[12][14][8] <= img[5264];\
        in_img_array[12][14][9] <= img[5265];\
        in_img_array[12][14][10] <= img[5266];\
        in_img_array[12][14][11] <= img[5267];\
        in_img_array[12][14][12] <= img[5268];\
        in_img_array[12][14][13] <= img[5269];\
        in_img_array[12][14][14] <= img[5270];\
        in_img_array[12][14][15] <= img[5271];\
        in_img_array[12][14][16] <= img[5272];\
        in_img_array[12][14][17] <= img[5273];\
        in_img_array[12][15][0] <= img[5274];\
        in_img_array[12][15][1] <= img[5275];\
        in_img_array[12][15][2] <= img[5276];\
        in_img_array[12][15][3] <= img[5277];\
        in_img_array[12][15][4] <= img[5278];\
        in_img_array[12][15][5] <= img[5279];\
        in_img_array[12][15][6] <= img[5280];\
        in_img_array[12][15][7] <= img[5281];\
        in_img_array[12][15][8] <= img[5282];\
        in_img_array[12][15][9] <= img[5283];\
        in_img_array[12][15][10] <= img[5284];\
        in_img_array[12][15][11] <= img[5285];\
        in_img_array[12][15][12] <= img[5286];\
        in_img_array[12][15][13] <= img[5287];\
        in_img_array[12][15][14] <= img[5288];\
        in_img_array[12][15][15] <= img[5289];\
        in_img_array[12][15][16] <= img[5290];\
        in_img_array[12][15][17] <= img[5291];\
        in_img_array[12][16][0] <= img[5292];\
        in_img_array[12][16][1] <= img[5293];\
        in_img_array[12][16][2] <= img[5294];\
        in_img_array[12][16][3] <= img[5295];\
        in_img_array[12][16][4] <= img[5296];\
        in_img_array[12][16][5] <= img[5297];\
        in_img_array[12][16][6] <= img[5298];\
        in_img_array[12][16][7] <= img[5299];\
        in_img_array[12][16][8] <= img[5300];\
        in_img_array[12][16][9] <= img[5301];\
        in_img_array[12][16][10] <= img[5302];\
        in_img_array[12][16][11] <= img[5303];\
        in_img_array[12][16][12] <= img[5304];\
        in_img_array[12][16][13] <= img[5305];\
        in_img_array[12][16][14] <= img[5306];\
        in_img_array[12][16][15] <= img[5307];\
        in_img_array[12][16][16] <= img[5308];\
        in_img_array[12][16][17] <= img[5309];\
        in_img_array[12][17][0] <= img[5310];\
        in_img_array[12][17][1] <= img[5311];\
        in_img_array[12][17][2] <= img[5312];\
        in_img_array[12][17][3] <= img[5313];\
        in_img_array[12][17][4] <= img[5314];\
        in_img_array[12][17][5] <= img[5315];\
        in_img_array[12][17][6] <= img[5316];\
        in_img_array[12][17][7] <= img[5317];\
        in_img_array[12][17][8] <= img[5318];\
        in_img_array[12][17][9] <= img[5319];\
        in_img_array[12][17][10] <= img[5320];\
        in_img_array[12][17][11] <= img[5321];\
        in_img_array[12][17][12] <= img[5322];\
        in_img_array[12][17][13] <= img[5323];\
        in_img_array[12][17][14] <= img[5324];\
        in_img_array[12][17][15] <= img[5325];\
        in_img_array[12][17][16] <= img[5326];\
        in_img_array[12][17][17] <= img[5327];\
        in_img_array[12][18][0] <= img[5328];\
        in_img_array[12][18][1] <= img[5329];\
        in_img_array[12][18][2] <= img[5330];\
        in_img_array[12][18][3] <= img[5331];\
        in_img_array[12][18][4] <= img[5332];\
        in_img_array[12][18][5] <= img[5333];\
        in_img_array[12][18][6] <= img[5334];\
        in_img_array[12][18][7] <= img[5335];\
        in_img_array[12][18][8] <= img[5336];\
        in_img_array[12][18][9] <= img[5337];\
        in_img_array[12][18][10] <= img[5338];\
        in_img_array[12][18][11] <= img[5339];\
        in_img_array[12][18][12] <= img[5340];\
        in_img_array[12][18][13] <= img[5341];\
        in_img_array[12][18][14] <= img[5342];\
        in_img_array[12][18][15] <= img[5343];\
        in_img_array[12][18][16] <= img[5344];\
        in_img_array[12][18][17] <= img[5345];\
        in_img_array[12][19][0] <= img[5346];\
        in_img_array[12][19][1] <= img[5347];\
        in_img_array[12][19][2] <= img[5348];\
        in_img_array[12][19][3] <= img[5349];\
        in_img_array[12][19][4] <= img[5350];\
        in_img_array[12][19][5] <= img[5351];\
        in_img_array[12][19][6] <= img[5352];\
        in_img_array[12][19][7] <= img[5353];\
        in_img_array[12][19][8] <= img[5354];\
        in_img_array[12][19][9] <= img[5355];\
        in_img_array[12][19][10] <= img[5356];\
        in_img_array[12][19][11] <= img[5357];\
        in_img_array[12][19][12] <= img[5358];\
        in_img_array[12][19][13] <= img[5359];\
        in_img_array[12][19][14] <= img[5360];\
        in_img_array[12][19][15] <= img[5361];\
        in_img_array[12][19][16] <= img[5362];\
        in_img_array[12][19][17] <= img[5363];\
        in_img_array[12][20][0] <= img[5364];\
        in_img_array[12][20][1] <= img[5365];\
        in_img_array[12][20][2] <= img[5366];\
        in_img_array[12][20][3] <= img[5367];\
        in_img_array[12][20][4] <= img[5368];\
        in_img_array[12][20][5] <= img[5369];\
        in_img_array[12][20][6] <= img[5370];\
        in_img_array[12][20][7] <= img[5371];\
        in_img_array[12][20][8] <= img[5372];\
        in_img_array[12][20][9] <= img[5373];\
        in_img_array[12][20][10] <= img[5374];\
        in_img_array[12][20][11] <= img[5375];\
        in_img_array[12][20][12] <= img[5376];\
        in_img_array[12][20][13] <= img[5377];\
        in_img_array[12][20][14] <= img[5378];\
        in_img_array[12][20][15] <= img[5379];\
        in_img_array[12][20][16] <= img[5380];\
        in_img_array[12][20][17] <= img[5381];\
        in_img_array[12][21][0] <= img[5382];\
        in_img_array[12][21][1] <= img[5383];\
        in_img_array[12][21][2] <= img[5384];\
        in_img_array[12][21][3] <= img[5385];\
        in_img_array[12][21][4] <= img[5386];\
        in_img_array[12][21][5] <= img[5387];\
        in_img_array[12][21][6] <= img[5388];\
        in_img_array[12][21][7] <= img[5389];\
        in_img_array[12][21][8] <= img[5390];\
        in_img_array[12][21][9] <= img[5391];\
        in_img_array[12][21][10] <= img[5392];\
        in_img_array[12][21][11] <= img[5393];\
        in_img_array[12][21][12] <= img[5394];\
        in_img_array[12][21][13] <= img[5395];\
        in_img_array[12][21][14] <= img[5396];\
        in_img_array[12][21][15] <= img[5397];\
        in_img_array[12][21][16] <= img[5398];\
        in_img_array[12][21][17] <= img[5399];\
        in_img_array[12][22][0] <= img[5400];\
        in_img_array[12][22][1] <= img[5401];\
        in_img_array[12][22][2] <= img[5402];\
        in_img_array[12][22][3] <= img[5403];\
        in_img_array[12][22][4] <= img[5404];\
        in_img_array[12][22][5] <= img[5405];\
        in_img_array[12][22][6] <= img[5406];\
        in_img_array[12][22][7] <= img[5407];\
        in_img_array[12][22][8] <= img[5408];\
        in_img_array[12][22][9] <= img[5409];\
        in_img_array[12][22][10] <= img[5410];\
        in_img_array[12][22][11] <= img[5411];\
        in_img_array[12][22][12] <= img[5412];\
        in_img_array[12][22][13] <= img[5413];\
        in_img_array[12][22][14] <= img[5414];\
        in_img_array[12][22][15] <= img[5415];\
        in_img_array[12][22][16] <= img[5416];\
        in_img_array[12][22][17] <= img[5417];\
        in_img_array[12][23][0] <= img[5418];\
        in_img_array[12][23][1] <= img[5419];\
        in_img_array[12][23][2] <= img[5420];\
        in_img_array[12][23][3] <= img[5421];\
        in_img_array[12][23][4] <= img[5422];\
        in_img_array[12][23][5] <= img[5423];\
        in_img_array[12][23][6] <= img[5424];\
        in_img_array[12][23][7] <= img[5425];\
        in_img_array[12][23][8] <= img[5426];\
        in_img_array[12][23][9] <= img[5427];\
        in_img_array[12][23][10] <= img[5428];\
        in_img_array[12][23][11] <= img[5429];\
        in_img_array[12][23][12] <= img[5430];\
        in_img_array[12][23][13] <= img[5431];\
        in_img_array[12][23][14] <= img[5432];\
        in_img_array[12][23][15] <= img[5433];\
        in_img_array[12][23][16] <= img[5434];\
        in_img_array[12][23][17] <= img[5435];\
        in_img_array[12][24][0] <= img[5436];\
        in_img_array[12][24][1] <= img[5437];\
        in_img_array[12][24][2] <= img[5438];\
        in_img_array[12][24][3] <= img[5439];\
        in_img_array[12][24][4] <= img[5440];\
        in_img_array[12][24][5] <= img[5441];\
        in_img_array[12][24][6] <= img[5442];\
        in_img_array[12][24][7] <= img[5443];\
        in_img_array[12][24][8] <= img[5444];\
        in_img_array[12][24][9] <= img[5445];\
        in_img_array[12][24][10] <= img[5446];\
        in_img_array[12][24][11] <= img[5447];\
        in_img_array[12][24][12] <= img[5448];\
        in_img_array[12][24][13] <= img[5449];\
        in_img_array[12][24][14] <= img[5450];\
        in_img_array[12][24][15] <= img[5451];\
        in_img_array[12][24][16] <= img[5452];\
        in_img_array[12][24][17] <= img[5453];\
        in_img_array[12][25][0] <= img[5454];\
        in_img_array[12][25][1] <= img[5455];\
        in_img_array[12][25][2] <= img[5456];\
        in_img_array[12][25][3] <= img[5457];\
        in_img_array[12][25][4] <= img[5458];\
        in_img_array[12][25][5] <= img[5459];\
        in_img_array[12][25][6] <= img[5460];\
        in_img_array[12][25][7] <= img[5461];\
        in_img_array[12][25][8] <= img[5462];\
        in_img_array[12][25][9] <= img[5463];\
        in_img_array[12][25][10] <= img[5464];\
        in_img_array[12][25][11] <= img[5465];\
        in_img_array[12][25][12] <= img[5466];\
        in_img_array[12][25][13] <= img[5467];\
        in_img_array[12][25][14] <= img[5468];\
        in_img_array[12][25][15] <= img[5469];\
        in_img_array[12][25][16] <= img[5470];\
        in_img_array[12][25][17] <= img[5471];\
        in_img_array[12][26][0] <= img[5472];\
        in_img_array[12][26][1] <= img[5473];\
        in_img_array[12][26][2] <= img[5474];\
        in_img_array[12][26][3] <= img[5475];\
        in_img_array[12][26][4] <= img[5476];\
        in_img_array[12][26][5] <= img[5477];\
        in_img_array[12][26][6] <= img[5478];\
        in_img_array[12][26][7] <= img[5479];\
        in_img_array[12][26][8] <= img[5480];\
        in_img_array[12][26][9] <= img[5481];\
        in_img_array[12][26][10] <= img[5482];\
        in_img_array[12][26][11] <= img[5483];\
        in_img_array[12][26][12] <= img[5484];\
        in_img_array[12][26][13] <= img[5485];\
        in_img_array[12][26][14] <= img[5486];\
        in_img_array[12][26][15] <= img[5487];\
        in_img_array[12][26][16] <= img[5488];\
        in_img_array[12][26][17] <= img[5489];\
        in_img_array[12][27][0] <= img[5490];\
        in_img_array[12][27][1] <= img[5491];\
        in_img_array[12][27][2] <= img[5492];\
        in_img_array[12][27][3] <= img[5493];\
        in_img_array[12][27][4] <= img[5494];\
        in_img_array[12][27][5] <= img[5495];\
        in_img_array[12][27][6] <= img[5496];\
        in_img_array[12][27][7] <= img[5497];\
        in_img_array[12][27][8] <= img[5498];\
        in_img_array[12][27][9] <= img[5499];\
        in_img_array[12][27][10] <= img[5500];\
        in_img_array[12][27][11] <= img[5501];\
        in_img_array[12][27][12] <= img[5502];\
        in_img_array[12][27][13] <= img[5503];\
        in_img_array[12][27][14] <= img[5504];\
        in_img_array[12][27][15] <= img[5505];\
        in_img_array[12][27][16] <= img[5506];\
        in_img_array[12][27][17] <= img[5507];\
        in_img_array[12][28][0] <= img[5508];\
        in_img_array[12][28][1] <= img[5509];\
        in_img_array[12][28][2] <= img[5510];\
        in_img_array[12][28][3] <= img[5511];\
        in_img_array[12][28][4] <= img[5512];\
        in_img_array[12][28][5] <= img[5513];\
        in_img_array[12][28][6] <= img[5514];\
        in_img_array[12][28][7] <= img[5515];\
        in_img_array[12][28][8] <= img[5516];\
        in_img_array[12][28][9] <= img[5517];\
        in_img_array[12][28][10] <= img[5518];\
        in_img_array[12][28][11] <= img[5519];\
        in_img_array[12][28][12] <= img[5520];\
        in_img_array[12][28][13] <= img[5521];\
        in_img_array[12][28][14] <= img[5522];\
        in_img_array[12][28][15] <= img[5523];\
        in_img_array[12][28][16] <= img[5524];\
        in_img_array[12][28][17] <= img[5525];\
        in_img_array[12][29][0] <= img[5526];\
        in_img_array[12][29][1] <= img[5527];\
        in_img_array[12][29][2] <= img[5528];\
        in_img_array[12][29][3] <= img[5529];\
        in_img_array[12][29][4] <= img[5530];\
        in_img_array[12][29][5] <= img[5531];\
        in_img_array[12][29][6] <= img[5532];\
        in_img_array[12][29][7] <= img[5533];\
        in_img_array[12][29][8] <= img[5534];\
        in_img_array[12][29][9] <= img[5535];\
        in_img_array[12][29][10] <= img[5536];\
        in_img_array[12][29][11] <= img[5537];\
        in_img_array[12][29][12] <= img[5538];\
        in_img_array[12][29][13] <= img[5539];\
        in_img_array[12][29][14] <= img[5540];\
        in_img_array[12][29][15] <= img[5541];\
        in_img_array[12][29][16] <= img[5542];\
        in_img_array[12][29][17] <= img[5543];\
        in_img_array[13][2][0] <= img[5544];\
        in_img_array[13][2][1] <= img[5545];\
        in_img_array[13][2][2] <= img[5546];\
        in_img_array[13][2][3] <= img[5547];\
        in_img_array[13][2][4] <= img[5548];\
        in_img_array[13][2][5] <= img[5549];\
        in_img_array[13][2][6] <= img[5550];\
        in_img_array[13][2][7] <= img[5551];\
        in_img_array[13][2][8] <= img[5552];\
        in_img_array[13][2][9] <= img[5553];\
        in_img_array[13][2][10] <= img[5554];\
        in_img_array[13][2][11] <= img[5555];\
        in_img_array[13][2][12] <= img[5556];\
        in_img_array[13][2][13] <= img[5557];\
        in_img_array[13][2][14] <= img[5558];\
        in_img_array[13][2][15] <= img[5559];\
        in_img_array[13][2][16] <= img[5560];\
        in_img_array[13][2][17] <= img[5561];\
        in_img_array[13][3][0] <= img[5562];\
        in_img_array[13][3][1] <= img[5563];\
        in_img_array[13][3][2] <= img[5564];\
        in_img_array[13][3][3] <= img[5565];\
        in_img_array[13][3][4] <= img[5566];\
        in_img_array[13][3][5] <= img[5567];\
        in_img_array[13][3][6] <= img[5568];\
        in_img_array[13][3][7] <= img[5569];\
        in_img_array[13][3][8] <= img[5570];\
        in_img_array[13][3][9] <= img[5571];\
        in_img_array[13][3][10] <= img[5572];\
        in_img_array[13][3][11] <= img[5573];\
        in_img_array[13][3][12] <= img[5574];\
        in_img_array[13][3][13] <= img[5575];\
        in_img_array[13][3][14] <= img[5576];\
        in_img_array[13][3][15] <= img[5577];\
        in_img_array[13][3][16] <= img[5578];\
        in_img_array[13][3][17] <= img[5579];\
        in_img_array[13][4][0] <= img[5580];\
        in_img_array[13][4][1] <= img[5581];\
        in_img_array[13][4][2] <= img[5582];\
        in_img_array[13][4][3] <= img[5583];\
        in_img_array[13][4][4] <= img[5584];\
        in_img_array[13][4][5] <= img[5585];\
        in_img_array[13][4][6] <= img[5586];\
        in_img_array[13][4][7] <= img[5587];\
        in_img_array[13][4][8] <= img[5588];\
        in_img_array[13][4][9] <= img[5589];\
        in_img_array[13][4][10] <= img[5590];\
        in_img_array[13][4][11] <= img[5591];\
        in_img_array[13][4][12] <= img[5592];\
        in_img_array[13][4][13] <= img[5593];\
        in_img_array[13][4][14] <= img[5594];\
        in_img_array[13][4][15] <= img[5595];\
        in_img_array[13][4][16] <= img[5596];\
        in_img_array[13][4][17] <= img[5597];\
        in_img_array[13][5][0] <= img[5598];\
        in_img_array[13][5][1] <= img[5599];\
        in_img_array[13][5][2] <= img[5600];\
        in_img_array[13][5][3] <= img[5601];\
        in_img_array[13][5][4] <= img[5602];\
        in_img_array[13][5][5] <= img[5603];\
        in_img_array[13][5][6] <= img[5604];\
        in_img_array[13][5][7] <= img[5605];\
        in_img_array[13][5][8] <= img[5606];\
        in_img_array[13][5][9] <= img[5607];\
        in_img_array[13][5][10] <= img[5608];\
        in_img_array[13][5][11] <= img[5609];\
        in_img_array[13][5][12] <= img[5610];\
        in_img_array[13][5][13] <= img[5611];\
        in_img_array[13][5][14] <= img[5612];\
        in_img_array[13][5][15] <= img[5613];\
        in_img_array[13][5][16] <= img[5614];\
        in_img_array[13][5][17] <= img[5615];\
        in_img_array[13][6][0] <= img[5616];\
        in_img_array[13][6][1] <= img[5617];\
        in_img_array[13][6][2] <= img[5618];\
        in_img_array[13][6][3] <= img[5619];\
        in_img_array[13][6][4] <= img[5620];\
        in_img_array[13][6][5] <= img[5621];\
        in_img_array[13][6][6] <= img[5622];\
        in_img_array[13][6][7] <= img[5623];\
        in_img_array[13][6][8] <= img[5624];\
        in_img_array[13][6][9] <= img[5625];\
        in_img_array[13][6][10] <= img[5626];\
        in_img_array[13][6][11] <= img[5627];\
        in_img_array[13][6][12] <= img[5628];\
        in_img_array[13][6][13] <= img[5629];\
        in_img_array[13][6][14] <= img[5630];\
        in_img_array[13][6][15] <= img[5631];\
        in_img_array[13][6][16] <= img[5632];\
        in_img_array[13][6][17] <= img[5633];\
        in_img_array[13][7][0] <= img[5634];\
        in_img_array[13][7][1] <= img[5635];\
        in_img_array[13][7][2] <= img[5636];\
        in_img_array[13][7][3] <= img[5637];\
        in_img_array[13][7][4] <= img[5638];\
        in_img_array[13][7][5] <= img[5639];\
        in_img_array[13][7][6] <= img[5640];\
        in_img_array[13][7][7] <= img[5641];\
        in_img_array[13][7][8] <= img[5642];\
        in_img_array[13][7][9] <= img[5643];\
        in_img_array[13][7][10] <= img[5644];\
        in_img_array[13][7][11] <= img[5645];\
        in_img_array[13][7][12] <= img[5646];\
        in_img_array[13][7][13] <= img[5647];\
        in_img_array[13][7][14] <= img[5648];\
        in_img_array[13][7][15] <= img[5649];\
        in_img_array[13][7][16] <= img[5650];\
        in_img_array[13][7][17] <= img[5651];\
        in_img_array[13][8][0] <= img[5652];\
        in_img_array[13][8][1] <= img[5653];\
        in_img_array[13][8][2] <= img[5654];\
        in_img_array[13][8][3] <= img[5655];\
        in_img_array[13][8][4] <= img[5656];\
        in_img_array[13][8][5] <= img[5657];\
        in_img_array[13][8][6] <= img[5658];\
        in_img_array[13][8][7] <= img[5659];\
        in_img_array[13][8][8] <= img[5660];\
        in_img_array[13][8][9] <= img[5661];\
        in_img_array[13][8][10] <= img[5662];\
        in_img_array[13][8][11] <= img[5663];\
        in_img_array[13][8][12] <= img[5664];\
        in_img_array[13][8][13] <= img[5665];\
        in_img_array[13][8][14] <= img[5666];\
        in_img_array[13][8][15] <= img[5667];\
        in_img_array[13][8][16] <= img[5668];\
        in_img_array[13][8][17] <= img[5669];\
        in_img_array[13][9][0] <= img[5670];\
        in_img_array[13][9][1] <= img[5671];\
        in_img_array[13][9][2] <= img[5672];\
        in_img_array[13][9][3] <= img[5673];\
        in_img_array[13][9][4] <= img[5674];\
        in_img_array[13][9][5] <= img[5675];\
        in_img_array[13][9][6] <= img[5676];\
        in_img_array[13][9][7] <= img[5677];\
        in_img_array[13][9][8] <= img[5678];\
        in_img_array[13][9][9] <= img[5679];\
        in_img_array[13][9][10] <= img[5680];\
        in_img_array[13][9][11] <= img[5681];\
        in_img_array[13][9][12] <= img[5682];\
        in_img_array[13][9][13] <= img[5683];\
        in_img_array[13][9][14] <= img[5684];\
        in_img_array[13][9][15] <= img[5685];\
        in_img_array[13][9][16] <= img[5686];\
        in_img_array[13][9][17] <= img[5687];\
        in_img_array[13][10][0] <= img[5688];\
        in_img_array[13][10][1] <= img[5689];\
        in_img_array[13][10][2] <= img[5690];\
        in_img_array[13][10][3] <= img[5691];\
        in_img_array[13][10][4] <= img[5692];\
        in_img_array[13][10][5] <= img[5693];\
        in_img_array[13][10][6] <= img[5694];\
        in_img_array[13][10][7] <= img[5695];\
        in_img_array[13][10][8] <= img[5696];\
        in_img_array[13][10][9] <= img[5697];\
        in_img_array[13][10][10] <= img[5698];\
        in_img_array[13][10][11] <= img[5699];\
        in_img_array[13][10][12] <= img[5700];\
        in_img_array[13][10][13] <= img[5701];\
        in_img_array[13][10][14] <= img[5702];\
        in_img_array[13][10][15] <= img[5703];\
        in_img_array[13][10][16] <= img[5704];\
        in_img_array[13][10][17] <= img[5705];\
        in_img_array[13][11][0] <= img[5706];\
        in_img_array[13][11][1] <= img[5707];\
        in_img_array[13][11][2] <= img[5708];\
        in_img_array[13][11][3] <= img[5709];\
        in_img_array[13][11][4] <= img[5710];\
        in_img_array[13][11][5] <= img[5711];\
        in_img_array[13][11][6] <= img[5712];\
        in_img_array[13][11][7] <= img[5713];\
        in_img_array[13][11][8] <= img[5714];\
        in_img_array[13][11][9] <= img[5715];\
        in_img_array[13][11][10] <= img[5716];\
        in_img_array[13][11][11] <= img[5717];\
        in_img_array[13][11][12] <= img[5718];\
        in_img_array[13][11][13] <= img[5719];\
        in_img_array[13][11][14] <= img[5720];\
        in_img_array[13][11][15] <= img[5721];\
        in_img_array[13][11][16] <= img[5722];\
        in_img_array[13][11][17] <= img[5723];\
        in_img_array[13][12][0] <= img[5724];\
        in_img_array[13][12][1] <= img[5725];\
        in_img_array[13][12][2] <= img[5726];\
        in_img_array[13][12][3] <= img[5727];\
        in_img_array[13][12][4] <= img[5728];\
        in_img_array[13][12][5] <= img[5729];\
        in_img_array[13][12][6] <= img[5730];\
        in_img_array[13][12][7] <= img[5731];\
        in_img_array[13][12][8] <= img[5732];\
        in_img_array[13][12][9] <= img[5733];\
        in_img_array[13][12][10] <= img[5734];\
        in_img_array[13][12][11] <= img[5735];\
        in_img_array[13][12][12] <= img[5736];\
        in_img_array[13][12][13] <= img[5737];\
        in_img_array[13][12][14] <= img[5738];\
        in_img_array[13][12][15] <= img[5739];\
        in_img_array[13][12][16] <= img[5740];\
        in_img_array[13][12][17] <= img[5741];\
        in_img_array[13][13][0] <= img[5742];\
        in_img_array[13][13][1] <= img[5743];\
        in_img_array[13][13][2] <= img[5744];\
        in_img_array[13][13][3] <= img[5745];\
        in_img_array[13][13][4] <= img[5746];\
        in_img_array[13][13][5] <= img[5747];\
        in_img_array[13][13][6] <= img[5748];\
        in_img_array[13][13][7] <= img[5749];\
        in_img_array[13][13][8] <= img[5750];\
        in_img_array[13][13][9] <= img[5751];\
        in_img_array[13][13][10] <= img[5752];\
        in_img_array[13][13][11] <= img[5753];\
        in_img_array[13][13][12] <= img[5754];\
        in_img_array[13][13][13] <= img[5755];\
        in_img_array[13][13][14] <= img[5756];\
        in_img_array[13][13][15] <= img[5757];\
        in_img_array[13][13][16] <= img[5758];\
        in_img_array[13][13][17] <= img[5759];\
        in_img_array[13][14][0] <= img[5760];\
        in_img_array[13][14][1] <= img[5761];\
        in_img_array[13][14][2] <= img[5762];\
        in_img_array[13][14][3] <= img[5763];\
        in_img_array[13][14][4] <= img[5764];\
        in_img_array[13][14][5] <= img[5765];\
        in_img_array[13][14][6] <= img[5766];\
        in_img_array[13][14][7] <= img[5767];\
        in_img_array[13][14][8] <= img[5768];\
        in_img_array[13][14][9] <= img[5769];\
        in_img_array[13][14][10] <= img[5770];\
        in_img_array[13][14][11] <= img[5771];\
        in_img_array[13][14][12] <= img[5772];\
        in_img_array[13][14][13] <= img[5773];\
        in_img_array[13][14][14] <= img[5774];\
        in_img_array[13][14][15] <= img[5775];\
        in_img_array[13][14][16] <= img[5776];\
        in_img_array[13][14][17] <= img[5777];\
        in_img_array[13][15][0] <= img[5778];\
        in_img_array[13][15][1] <= img[5779];\
        in_img_array[13][15][2] <= img[5780];\
        in_img_array[13][15][3] <= img[5781];\
        in_img_array[13][15][4] <= img[5782];\
        in_img_array[13][15][5] <= img[5783];\
        in_img_array[13][15][6] <= img[5784];\
        in_img_array[13][15][7] <= img[5785];\
        in_img_array[13][15][8] <= img[5786];\
        in_img_array[13][15][9] <= img[5787];\
        in_img_array[13][15][10] <= img[5788];\
        in_img_array[13][15][11] <= img[5789];\
        in_img_array[13][15][12] <= img[5790];\
        in_img_array[13][15][13] <= img[5791];\
        in_img_array[13][15][14] <= img[5792];\
        in_img_array[13][15][15] <= img[5793];\
        in_img_array[13][15][16] <= img[5794];\
        in_img_array[13][15][17] <= img[5795];\
        in_img_array[13][16][0] <= img[5796];\
        in_img_array[13][16][1] <= img[5797];\
        in_img_array[13][16][2] <= img[5798];\
        in_img_array[13][16][3] <= img[5799];\
        in_img_array[13][16][4] <= img[5800];\
        in_img_array[13][16][5] <= img[5801];\
        in_img_array[13][16][6] <= img[5802];\
        in_img_array[13][16][7] <= img[5803];\
        in_img_array[13][16][8] <= img[5804];\
        in_img_array[13][16][9] <= img[5805];\
        in_img_array[13][16][10] <= img[5806];\
        in_img_array[13][16][11] <= img[5807];\
        in_img_array[13][16][12] <= img[5808];\
        in_img_array[13][16][13] <= img[5809];\
        in_img_array[13][16][14] <= img[5810];\
        in_img_array[13][16][15] <= img[5811];\
        in_img_array[13][16][16] <= img[5812];\
        in_img_array[13][16][17] <= img[5813];\
        in_img_array[13][17][0] <= img[5814];\
        in_img_array[13][17][1] <= img[5815];\
        in_img_array[13][17][2] <= img[5816];\
        in_img_array[13][17][3] <= img[5817];\
        in_img_array[13][17][4] <= img[5818];\
        in_img_array[13][17][5] <= img[5819];\
        in_img_array[13][17][6] <= img[5820];\
        in_img_array[13][17][7] <= img[5821];\
        in_img_array[13][17][8] <= img[5822];\
        in_img_array[13][17][9] <= img[5823];\
        in_img_array[13][17][10] <= img[5824];\
        in_img_array[13][17][11] <= img[5825];\
        in_img_array[13][17][12] <= img[5826];\
        in_img_array[13][17][13] <= img[5827];\
        in_img_array[13][17][14] <= img[5828];\
        in_img_array[13][17][15] <= img[5829];\
        in_img_array[13][17][16] <= img[5830];\
        in_img_array[13][17][17] <= img[5831];\
        in_img_array[13][18][0] <= img[5832];\
        in_img_array[13][18][1] <= img[5833];\
        in_img_array[13][18][2] <= img[5834];\
        in_img_array[13][18][3] <= img[5835];\
        in_img_array[13][18][4] <= img[5836];\
        in_img_array[13][18][5] <= img[5837];\
        in_img_array[13][18][6] <= img[5838];\
        in_img_array[13][18][7] <= img[5839];\
        in_img_array[13][18][8] <= img[5840];\
        in_img_array[13][18][9] <= img[5841];\
        in_img_array[13][18][10] <= img[5842];\
        in_img_array[13][18][11] <= img[5843];\
        in_img_array[13][18][12] <= img[5844];\
        in_img_array[13][18][13] <= img[5845];\
        in_img_array[13][18][14] <= img[5846];\
        in_img_array[13][18][15] <= img[5847];\
        in_img_array[13][18][16] <= img[5848];\
        in_img_array[13][18][17] <= img[5849];\
        in_img_array[13][19][0] <= img[5850];\
        in_img_array[13][19][1] <= img[5851];\
        in_img_array[13][19][2] <= img[5852];\
        in_img_array[13][19][3] <= img[5853];\
        in_img_array[13][19][4] <= img[5854];\
        in_img_array[13][19][5] <= img[5855];\
        in_img_array[13][19][6] <= img[5856];\
        in_img_array[13][19][7] <= img[5857];\
        in_img_array[13][19][8] <= img[5858];\
        in_img_array[13][19][9] <= img[5859];\
        in_img_array[13][19][10] <= img[5860];\
        in_img_array[13][19][11] <= img[5861];\
        in_img_array[13][19][12] <= img[5862];\
        in_img_array[13][19][13] <= img[5863];\
        in_img_array[13][19][14] <= img[5864];\
        in_img_array[13][19][15] <= img[5865];\
        in_img_array[13][19][16] <= img[5866];\
        in_img_array[13][19][17] <= img[5867];\
        in_img_array[13][20][0] <= img[5868];\
        in_img_array[13][20][1] <= img[5869];\
        in_img_array[13][20][2] <= img[5870];\
        in_img_array[13][20][3] <= img[5871];\
        in_img_array[13][20][4] <= img[5872];\
        in_img_array[13][20][5] <= img[5873];\
        in_img_array[13][20][6] <= img[5874];\
        in_img_array[13][20][7] <= img[5875];\
        in_img_array[13][20][8] <= img[5876];\
        in_img_array[13][20][9] <= img[5877];\
        in_img_array[13][20][10] <= img[5878];\
        in_img_array[13][20][11] <= img[5879];\
        in_img_array[13][20][12] <= img[5880];\
        in_img_array[13][20][13] <= img[5881];\
        in_img_array[13][20][14] <= img[5882];\
        in_img_array[13][20][15] <= img[5883];\
        in_img_array[13][20][16] <= img[5884];\
        in_img_array[13][20][17] <= img[5885];\
        in_img_array[13][21][0] <= img[5886];\
        in_img_array[13][21][1] <= img[5887];\
        in_img_array[13][21][2] <= img[5888];\
        in_img_array[13][21][3] <= img[5889];\
        in_img_array[13][21][4] <= img[5890];\
        in_img_array[13][21][5] <= img[5891];\
        in_img_array[13][21][6] <= img[5892];\
        in_img_array[13][21][7] <= img[5893];\
        in_img_array[13][21][8] <= img[5894];\
        in_img_array[13][21][9] <= img[5895];\
        in_img_array[13][21][10] <= img[5896];\
        in_img_array[13][21][11] <= img[5897];\
        in_img_array[13][21][12] <= img[5898];\
        in_img_array[13][21][13] <= img[5899];\
        in_img_array[13][21][14] <= img[5900];\
        in_img_array[13][21][15] <= img[5901];\
        in_img_array[13][21][16] <= img[5902];\
        in_img_array[13][21][17] <= img[5903];\
        in_img_array[13][22][0] <= img[5904];\
        in_img_array[13][22][1] <= img[5905];\
        in_img_array[13][22][2] <= img[5906];\
        in_img_array[13][22][3] <= img[5907];\
        in_img_array[13][22][4] <= img[5908];\
        in_img_array[13][22][5] <= img[5909];\
        in_img_array[13][22][6] <= img[5910];\
        in_img_array[13][22][7] <= img[5911];\
        in_img_array[13][22][8] <= img[5912];\
        in_img_array[13][22][9] <= img[5913];\
        in_img_array[13][22][10] <= img[5914];\
        in_img_array[13][22][11] <= img[5915];\
        in_img_array[13][22][12] <= img[5916];\
        in_img_array[13][22][13] <= img[5917];\
        in_img_array[13][22][14] <= img[5918];\
        in_img_array[13][22][15] <= img[5919];\
        in_img_array[13][22][16] <= img[5920];\
        in_img_array[13][22][17] <= img[5921];\
        in_img_array[13][23][0] <= img[5922];\
        in_img_array[13][23][1] <= img[5923];\
        in_img_array[13][23][2] <= img[5924];\
        in_img_array[13][23][3] <= img[5925];\
        in_img_array[13][23][4] <= img[5926];\
        in_img_array[13][23][5] <= img[5927];\
        in_img_array[13][23][6] <= img[5928];\
        in_img_array[13][23][7] <= img[5929];\
        in_img_array[13][23][8] <= img[5930];\
        in_img_array[13][23][9] <= img[5931];\
        in_img_array[13][23][10] <= img[5932];\
        in_img_array[13][23][11] <= img[5933];\
        in_img_array[13][23][12] <= img[5934];\
        in_img_array[13][23][13] <= img[5935];\
        in_img_array[13][23][14] <= img[5936];\
        in_img_array[13][23][15] <= img[5937];\
        in_img_array[13][23][16] <= img[5938];\
        in_img_array[13][23][17] <= img[5939];\
        in_img_array[13][24][0] <= img[5940];\
        in_img_array[13][24][1] <= img[5941];\
        in_img_array[13][24][2] <= img[5942];\
        in_img_array[13][24][3] <= img[5943];\
        in_img_array[13][24][4] <= img[5944];\
        in_img_array[13][24][5] <= img[5945];\
        in_img_array[13][24][6] <= img[5946];\
        in_img_array[13][24][7] <= img[5947];\
        in_img_array[13][24][8] <= img[5948];\
        in_img_array[13][24][9] <= img[5949];\
        in_img_array[13][24][10] <= img[5950];\
        in_img_array[13][24][11] <= img[5951];\
        in_img_array[13][24][12] <= img[5952];\
        in_img_array[13][24][13] <= img[5953];\
        in_img_array[13][24][14] <= img[5954];\
        in_img_array[13][24][15] <= img[5955];\
        in_img_array[13][24][16] <= img[5956];\
        in_img_array[13][24][17] <= img[5957];\
        in_img_array[13][25][0] <= img[5958];\
        in_img_array[13][25][1] <= img[5959];\
        in_img_array[13][25][2] <= img[5960];\
        in_img_array[13][25][3] <= img[5961];\
        in_img_array[13][25][4] <= img[5962];\
        in_img_array[13][25][5] <= img[5963];\
        in_img_array[13][25][6] <= img[5964];\
        in_img_array[13][25][7] <= img[5965];\
        in_img_array[13][25][8] <= img[5966];\
        in_img_array[13][25][9] <= img[5967];\
        in_img_array[13][25][10] <= img[5968];\
        in_img_array[13][25][11] <= img[5969];\
        in_img_array[13][25][12] <= img[5970];\
        in_img_array[13][25][13] <= img[5971];\
        in_img_array[13][25][14] <= img[5972];\
        in_img_array[13][25][15] <= img[5973];\
        in_img_array[13][25][16] <= img[5974];\
        in_img_array[13][25][17] <= img[5975];\
        in_img_array[13][26][0] <= img[5976];\
        in_img_array[13][26][1] <= img[5977];\
        in_img_array[13][26][2] <= img[5978];\
        in_img_array[13][26][3] <= img[5979];\
        in_img_array[13][26][4] <= img[5980];\
        in_img_array[13][26][5] <= img[5981];\
        in_img_array[13][26][6] <= img[5982];\
        in_img_array[13][26][7] <= img[5983];\
        in_img_array[13][26][8] <= img[5984];\
        in_img_array[13][26][9] <= img[5985];\
        in_img_array[13][26][10] <= img[5986];\
        in_img_array[13][26][11] <= img[5987];\
        in_img_array[13][26][12] <= img[5988];\
        in_img_array[13][26][13] <= img[5989];\
        in_img_array[13][26][14] <= img[5990];\
        in_img_array[13][26][15] <= img[5991];\
        in_img_array[13][26][16] <= img[5992];\
        in_img_array[13][26][17] <= img[5993];\
        in_img_array[13][27][0] <= img[5994];\
        in_img_array[13][27][1] <= img[5995];\
        in_img_array[13][27][2] <= img[5996];\
        in_img_array[13][27][3] <= img[5997];\
        in_img_array[13][27][4] <= img[5998];\
        in_img_array[13][27][5] <= img[5999];\
        in_img_array[13][27][6] <= img[6000];\
        in_img_array[13][27][7] <= img[6001];\
        in_img_array[13][27][8] <= img[6002];\
        in_img_array[13][27][9] <= img[6003];\
        in_img_array[13][27][10] <= img[6004];\
        in_img_array[13][27][11] <= img[6005];\
        in_img_array[13][27][12] <= img[6006];\
        in_img_array[13][27][13] <= img[6007];\
        in_img_array[13][27][14] <= img[6008];\
        in_img_array[13][27][15] <= img[6009];\
        in_img_array[13][27][16] <= img[6010];\
        in_img_array[13][27][17] <= img[6011];\
        in_img_array[13][28][0] <= img[6012];\
        in_img_array[13][28][1] <= img[6013];\
        in_img_array[13][28][2] <= img[6014];\
        in_img_array[13][28][3] <= img[6015];\
        in_img_array[13][28][4] <= img[6016];\
        in_img_array[13][28][5] <= img[6017];\
        in_img_array[13][28][6] <= img[6018];\
        in_img_array[13][28][7] <= img[6019];\
        in_img_array[13][28][8] <= img[6020];\
        in_img_array[13][28][9] <= img[6021];\
        in_img_array[13][28][10] <= img[6022];\
        in_img_array[13][28][11] <= img[6023];\
        in_img_array[13][28][12] <= img[6024];\
        in_img_array[13][28][13] <= img[6025];\
        in_img_array[13][28][14] <= img[6026];\
        in_img_array[13][28][15] <= img[6027];\
        in_img_array[13][28][16] <= img[6028];\
        in_img_array[13][28][17] <= img[6029];\
        in_img_array[13][29][0] <= img[6030];\
        in_img_array[13][29][1] <= img[6031];\
        in_img_array[13][29][2] <= img[6032];\
        in_img_array[13][29][3] <= img[6033];\
        in_img_array[13][29][4] <= img[6034];\
        in_img_array[13][29][5] <= img[6035];\
        in_img_array[13][29][6] <= img[6036];\
        in_img_array[13][29][7] <= img[6037];\
        in_img_array[13][29][8] <= img[6038];\
        in_img_array[13][29][9] <= img[6039];\
        in_img_array[13][29][10] <= img[6040];\
        in_img_array[13][29][11] <= img[6041];\
        in_img_array[13][29][12] <= img[6042];\
        in_img_array[13][29][13] <= img[6043];\
        in_img_array[13][29][14] <= img[6044];\
        in_img_array[13][29][15] <= img[6045];\
        in_img_array[13][29][16] <= img[6046];\
        in_img_array[13][29][17] <= img[6047];\
        in_img_array[14][2][0] <= img[6048];\
        in_img_array[14][2][1] <= img[6049];\
        in_img_array[14][2][2] <= img[6050];\
        in_img_array[14][2][3] <= img[6051];\
        in_img_array[14][2][4] <= img[6052];\
        in_img_array[14][2][5] <= img[6053];\
        in_img_array[14][2][6] <= img[6054];\
        in_img_array[14][2][7] <= img[6055];\
        in_img_array[14][2][8] <= img[6056];\
        in_img_array[14][2][9] <= img[6057];\
        in_img_array[14][2][10] <= img[6058];\
        in_img_array[14][2][11] <= img[6059];\
        in_img_array[14][2][12] <= img[6060];\
        in_img_array[14][2][13] <= img[6061];\
        in_img_array[14][2][14] <= img[6062];\
        in_img_array[14][2][15] <= img[6063];\
        in_img_array[14][2][16] <= img[6064];\
        in_img_array[14][2][17] <= img[6065];\
        in_img_array[14][3][0] <= img[6066];\
        in_img_array[14][3][1] <= img[6067];\
        in_img_array[14][3][2] <= img[6068];\
        in_img_array[14][3][3] <= img[6069];\
        in_img_array[14][3][4] <= img[6070];\
        in_img_array[14][3][5] <= img[6071];\
        in_img_array[14][3][6] <= img[6072];\
        in_img_array[14][3][7] <= img[6073];\
        in_img_array[14][3][8] <= img[6074];\
        in_img_array[14][3][9] <= img[6075];\
        in_img_array[14][3][10] <= img[6076];\
        in_img_array[14][3][11] <= img[6077];\
        in_img_array[14][3][12] <= img[6078];\
        in_img_array[14][3][13] <= img[6079];\
        in_img_array[14][3][14] <= img[6080];\
        in_img_array[14][3][15] <= img[6081];\
        in_img_array[14][3][16] <= img[6082];\
        in_img_array[14][3][17] <= img[6083];\
        in_img_array[14][4][0] <= img[6084];\
        in_img_array[14][4][1] <= img[6085];\
        in_img_array[14][4][2] <= img[6086];\
        in_img_array[14][4][3] <= img[6087];\
        in_img_array[14][4][4] <= img[6088];\
        in_img_array[14][4][5] <= img[6089];\
        in_img_array[14][4][6] <= img[6090];\
        in_img_array[14][4][7] <= img[6091];\
        in_img_array[14][4][8] <= img[6092];\
        in_img_array[14][4][9] <= img[6093];\
        in_img_array[14][4][10] <= img[6094];\
        in_img_array[14][4][11] <= img[6095];\
        in_img_array[14][4][12] <= img[6096];\
        in_img_array[14][4][13] <= img[6097];\
        in_img_array[14][4][14] <= img[6098];\
        in_img_array[14][4][15] <= img[6099];\
        in_img_array[14][4][16] <= img[6100];\
        in_img_array[14][4][17] <= img[6101];\
        in_img_array[14][5][0] <= img[6102];\
        in_img_array[14][5][1] <= img[6103];\
        in_img_array[14][5][2] <= img[6104];\
        in_img_array[14][5][3] <= img[6105];\
        in_img_array[14][5][4] <= img[6106];\
        in_img_array[14][5][5] <= img[6107];\
        in_img_array[14][5][6] <= img[6108];\
        in_img_array[14][5][7] <= img[6109];\
        in_img_array[14][5][8] <= img[6110];\
        in_img_array[14][5][9] <= img[6111];\
        in_img_array[14][5][10] <= img[6112];\
        in_img_array[14][5][11] <= img[6113];\
        in_img_array[14][5][12] <= img[6114];\
        in_img_array[14][5][13] <= img[6115];\
        in_img_array[14][5][14] <= img[6116];\
        in_img_array[14][5][15] <= img[6117];\
        in_img_array[14][5][16] <= img[6118];\
        in_img_array[14][5][17] <= img[6119];\
        in_img_array[14][6][0] <= img[6120];\
        in_img_array[14][6][1] <= img[6121];\
        in_img_array[14][6][2] <= img[6122];\
        in_img_array[14][6][3] <= img[6123];\
        in_img_array[14][6][4] <= img[6124];\
        in_img_array[14][6][5] <= img[6125];\
        in_img_array[14][6][6] <= img[6126];\
        in_img_array[14][6][7] <= img[6127];\
        in_img_array[14][6][8] <= img[6128];\
        in_img_array[14][6][9] <= img[6129];\
        in_img_array[14][6][10] <= img[6130];\
        in_img_array[14][6][11] <= img[6131];\
        in_img_array[14][6][12] <= img[6132];\
        in_img_array[14][6][13] <= img[6133];\
        in_img_array[14][6][14] <= img[6134];\
        in_img_array[14][6][15] <= img[6135];\
        in_img_array[14][6][16] <= img[6136];\
        in_img_array[14][6][17] <= img[6137];\
        in_img_array[14][7][0] <= img[6138];\
        in_img_array[14][7][1] <= img[6139];\
        in_img_array[14][7][2] <= img[6140];\
        in_img_array[14][7][3] <= img[6141];\
        in_img_array[14][7][4] <= img[6142];\
        in_img_array[14][7][5] <= img[6143];\
        in_img_array[14][7][6] <= img[6144];\
        in_img_array[14][7][7] <= img[6145];\
        in_img_array[14][7][8] <= img[6146];\
        in_img_array[14][7][9] <= img[6147];\
        in_img_array[14][7][10] <= img[6148];\
        in_img_array[14][7][11] <= img[6149];\
        in_img_array[14][7][12] <= img[6150];\
        in_img_array[14][7][13] <= img[6151];\
        in_img_array[14][7][14] <= img[6152];\
        in_img_array[14][7][15] <= img[6153];\
        in_img_array[14][7][16] <= img[6154];\
        in_img_array[14][7][17] <= img[6155];\
        in_img_array[14][8][0] <= img[6156];\
        in_img_array[14][8][1] <= img[6157];\
        in_img_array[14][8][2] <= img[6158];\
        in_img_array[14][8][3] <= img[6159];\
        in_img_array[14][8][4] <= img[6160];\
        in_img_array[14][8][5] <= img[6161];\
        in_img_array[14][8][6] <= img[6162];\
        in_img_array[14][8][7] <= img[6163];\
        in_img_array[14][8][8] <= img[6164];\
        in_img_array[14][8][9] <= img[6165];\
        in_img_array[14][8][10] <= img[6166];\
        in_img_array[14][8][11] <= img[6167];\
        in_img_array[14][8][12] <= img[6168];\
        in_img_array[14][8][13] <= img[6169];\
        in_img_array[14][8][14] <= img[6170];\
        in_img_array[14][8][15] <= img[6171];\
        in_img_array[14][8][16] <= img[6172];\
        in_img_array[14][8][17] <= img[6173];\
        in_img_array[14][9][0] <= img[6174];\
        in_img_array[14][9][1] <= img[6175];\
        in_img_array[14][9][2] <= img[6176];\
        in_img_array[14][9][3] <= img[6177];\
        in_img_array[14][9][4] <= img[6178];\
        in_img_array[14][9][5] <= img[6179];\
        in_img_array[14][9][6] <= img[6180];\
        in_img_array[14][9][7] <= img[6181];\
        in_img_array[14][9][8] <= img[6182];\
        in_img_array[14][9][9] <= img[6183];\
        in_img_array[14][9][10] <= img[6184];\
        in_img_array[14][9][11] <= img[6185];\
        in_img_array[14][9][12] <= img[6186];\
        in_img_array[14][9][13] <= img[6187];\
        in_img_array[14][9][14] <= img[6188];\
        in_img_array[14][9][15] <= img[6189];\
        in_img_array[14][9][16] <= img[6190];\
        in_img_array[14][9][17] <= img[6191];\
        in_img_array[14][10][0] <= img[6192];\
        in_img_array[14][10][1] <= img[6193];\
        in_img_array[14][10][2] <= img[6194];\
        in_img_array[14][10][3] <= img[6195];\
        in_img_array[14][10][4] <= img[6196];\
        in_img_array[14][10][5] <= img[6197];\
        in_img_array[14][10][6] <= img[6198];\
        in_img_array[14][10][7] <= img[6199];\
        in_img_array[14][10][8] <= img[6200];\
        in_img_array[14][10][9] <= img[6201];\
        in_img_array[14][10][10] <= img[6202];\
        in_img_array[14][10][11] <= img[6203];\
        in_img_array[14][10][12] <= img[6204];\
        in_img_array[14][10][13] <= img[6205];\
        in_img_array[14][10][14] <= img[6206];\
        in_img_array[14][10][15] <= img[6207];\
        in_img_array[14][10][16] <= img[6208];\
        in_img_array[14][10][17] <= img[6209];\
        in_img_array[14][11][0] <= img[6210];\
        in_img_array[14][11][1] <= img[6211];\
        in_img_array[14][11][2] <= img[6212];\
        in_img_array[14][11][3] <= img[6213];\
        in_img_array[14][11][4] <= img[6214];\
        in_img_array[14][11][5] <= img[6215];\
        in_img_array[14][11][6] <= img[6216];\
        in_img_array[14][11][7] <= img[6217];\
        in_img_array[14][11][8] <= img[6218];\
        in_img_array[14][11][9] <= img[6219];\
        in_img_array[14][11][10] <= img[6220];\
        in_img_array[14][11][11] <= img[6221];\
        in_img_array[14][11][12] <= img[6222];\
        in_img_array[14][11][13] <= img[6223];\
        in_img_array[14][11][14] <= img[6224];\
        in_img_array[14][11][15] <= img[6225];\
        in_img_array[14][11][16] <= img[6226];\
        in_img_array[14][11][17] <= img[6227];\
        in_img_array[14][12][0] <= img[6228];\
        in_img_array[14][12][1] <= img[6229];\
        in_img_array[14][12][2] <= img[6230];\
        in_img_array[14][12][3] <= img[6231];\
        in_img_array[14][12][4] <= img[6232];\
        in_img_array[14][12][5] <= img[6233];\
        in_img_array[14][12][6] <= img[6234];\
        in_img_array[14][12][7] <= img[6235];\
        in_img_array[14][12][8] <= img[6236];\
        in_img_array[14][12][9] <= img[6237];\
        in_img_array[14][12][10] <= img[6238];\
        in_img_array[14][12][11] <= img[6239];\
        in_img_array[14][12][12] <= img[6240];\
        in_img_array[14][12][13] <= img[6241];\
        in_img_array[14][12][14] <= img[6242];\
        in_img_array[14][12][15] <= img[6243];\
        in_img_array[14][12][16] <= img[6244];\
        in_img_array[14][12][17] <= img[6245];\
        in_img_array[14][13][0] <= img[6246];\
        in_img_array[14][13][1] <= img[6247];\
        in_img_array[14][13][2] <= img[6248];\
        in_img_array[14][13][3] <= img[6249];\
        in_img_array[14][13][4] <= img[6250];\
        in_img_array[14][13][5] <= img[6251];\
        in_img_array[14][13][6] <= img[6252];\
        in_img_array[14][13][7] <= img[6253];\
        in_img_array[14][13][8] <= img[6254];\
        in_img_array[14][13][9] <= img[6255];\
        in_img_array[14][13][10] <= img[6256];\
        in_img_array[14][13][11] <= img[6257];\
        in_img_array[14][13][12] <= img[6258];\
        in_img_array[14][13][13] <= img[6259];\
        in_img_array[14][13][14] <= img[6260];\
        in_img_array[14][13][15] <= img[6261];\
        in_img_array[14][13][16] <= img[6262];\
        in_img_array[14][13][17] <= img[6263];\
        in_img_array[14][14][0] <= img[6264];\
        in_img_array[14][14][1] <= img[6265];\
        in_img_array[14][14][2] <= img[6266];\
        in_img_array[14][14][3] <= img[6267];\
        in_img_array[14][14][4] <= img[6268];\
        in_img_array[14][14][5] <= img[6269];\
        in_img_array[14][14][6] <= img[6270];\
        in_img_array[14][14][7] <= img[6271];\
        in_img_array[14][14][8] <= img[6272];\
        in_img_array[14][14][9] <= img[6273];\
        in_img_array[14][14][10] <= img[6274];\
        in_img_array[14][14][11] <= img[6275];\
        in_img_array[14][14][12] <= img[6276];\
        in_img_array[14][14][13] <= img[6277];\
        in_img_array[14][14][14] <= img[6278];\
        in_img_array[14][14][15] <= img[6279];\
        in_img_array[14][14][16] <= img[6280];\
        in_img_array[14][14][17] <= img[6281];\
        in_img_array[14][15][0] <= img[6282];\
        in_img_array[14][15][1] <= img[6283];\
        in_img_array[14][15][2] <= img[6284];\
        in_img_array[14][15][3] <= img[6285];\
        in_img_array[14][15][4] <= img[6286];\
        in_img_array[14][15][5] <= img[6287];\
        in_img_array[14][15][6] <= img[6288];\
        in_img_array[14][15][7] <= img[6289];\
        in_img_array[14][15][8] <= img[6290];\
        in_img_array[14][15][9] <= img[6291];\
        in_img_array[14][15][10] <= img[6292];\
        in_img_array[14][15][11] <= img[6293];\
        in_img_array[14][15][12] <= img[6294];\
        in_img_array[14][15][13] <= img[6295];\
        in_img_array[14][15][14] <= img[6296];\
        in_img_array[14][15][15] <= img[6297];\
        in_img_array[14][15][16] <= img[6298];\
        in_img_array[14][15][17] <= img[6299];\
        in_img_array[14][16][0] <= img[6300];\
        in_img_array[14][16][1] <= img[6301];\
        in_img_array[14][16][2] <= img[6302];\
        in_img_array[14][16][3] <= img[6303];\
        in_img_array[14][16][4] <= img[6304];\
        in_img_array[14][16][5] <= img[6305];\
        in_img_array[14][16][6] <= img[6306];\
        in_img_array[14][16][7] <= img[6307];\
        in_img_array[14][16][8] <= img[6308];\
        in_img_array[14][16][9] <= img[6309];\
        in_img_array[14][16][10] <= img[6310];\
        in_img_array[14][16][11] <= img[6311];\
        in_img_array[14][16][12] <= img[6312];\
        in_img_array[14][16][13] <= img[6313];\
        in_img_array[14][16][14] <= img[6314];\
        in_img_array[14][16][15] <= img[6315];\
        in_img_array[14][16][16] <= img[6316];\
        in_img_array[14][16][17] <= img[6317];\
        in_img_array[14][17][0] <= img[6318];\
        in_img_array[14][17][1] <= img[6319];\
        in_img_array[14][17][2] <= img[6320];\
        in_img_array[14][17][3] <= img[6321];\
        in_img_array[14][17][4] <= img[6322];\
        in_img_array[14][17][5] <= img[6323];\
        in_img_array[14][17][6] <= img[6324];\
        in_img_array[14][17][7] <= img[6325];\
        in_img_array[14][17][8] <= img[6326];\
        in_img_array[14][17][9] <= img[6327];\
        in_img_array[14][17][10] <= img[6328];\
        in_img_array[14][17][11] <= img[6329];\
        in_img_array[14][17][12] <= img[6330];\
        in_img_array[14][17][13] <= img[6331];\
        in_img_array[14][17][14] <= img[6332];\
        in_img_array[14][17][15] <= img[6333];\
        in_img_array[14][17][16] <= img[6334];\
        in_img_array[14][17][17] <= img[6335];\
        in_img_array[14][18][0] <= img[6336];\
        in_img_array[14][18][1] <= img[6337];\
        in_img_array[14][18][2] <= img[6338];\
        in_img_array[14][18][3] <= img[6339];\
        in_img_array[14][18][4] <= img[6340];\
        in_img_array[14][18][5] <= img[6341];\
        in_img_array[14][18][6] <= img[6342];\
        in_img_array[14][18][7] <= img[6343];\
        in_img_array[14][18][8] <= img[6344];\
        in_img_array[14][18][9] <= img[6345];\
        in_img_array[14][18][10] <= img[6346];\
        in_img_array[14][18][11] <= img[6347];\
        in_img_array[14][18][12] <= img[6348];\
        in_img_array[14][18][13] <= img[6349];\
        in_img_array[14][18][14] <= img[6350];\
        in_img_array[14][18][15] <= img[6351];\
        in_img_array[14][18][16] <= img[6352];\
        in_img_array[14][18][17] <= img[6353];\
        in_img_array[14][19][0] <= img[6354];\
        in_img_array[14][19][1] <= img[6355];\
        in_img_array[14][19][2] <= img[6356];\
        in_img_array[14][19][3] <= img[6357];\
        in_img_array[14][19][4] <= img[6358];\
        in_img_array[14][19][5] <= img[6359];\
        in_img_array[14][19][6] <= img[6360];\
        in_img_array[14][19][7] <= img[6361];\
        in_img_array[14][19][8] <= img[6362];\
        in_img_array[14][19][9] <= img[6363];\
        in_img_array[14][19][10] <= img[6364];\
        in_img_array[14][19][11] <= img[6365];\
        in_img_array[14][19][12] <= img[6366];\
        in_img_array[14][19][13] <= img[6367];\
        in_img_array[14][19][14] <= img[6368];\
        in_img_array[14][19][15] <= img[6369];\
        in_img_array[14][19][16] <= img[6370];\
        in_img_array[14][19][17] <= img[6371];\
        in_img_array[14][20][0] <= img[6372];\
        in_img_array[14][20][1] <= img[6373];\
        in_img_array[14][20][2] <= img[6374];\
        in_img_array[14][20][3] <= img[6375];\
        in_img_array[14][20][4] <= img[6376];\
        in_img_array[14][20][5] <= img[6377];\
        in_img_array[14][20][6] <= img[6378];\
        in_img_array[14][20][7] <= img[6379];\
        in_img_array[14][20][8] <= img[6380];\
        in_img_array[14][20][9] <= img[6381];\
        in_img_array[14][20][10] <= img[6382];\
        in_img_array[14][20][11] <= img[6383];\
        in_img_array[14][20][12] <= img[6384];\
        in_img_array[14][20][13] <= img[6385];\
        in_img_array[14][20][14] <= img[6386];\
        in_img_array[14][20][15] <= img[6387];\
        in_img_array[14][20][16] <= img[6388];\
        in_img_array[14][20][17] <= img[6389];\
        in_img_array[14][21][0] <= img[6390];\
        in_img_array[14][21][1] <= img[6391];\
        in_img_array[14][21][2] <= img[6392];\
        in_img_array[14][21][3] <= img[6393];\
        in_img_array[14][21][4] <= img[6394];\
        in_img_array[14][21][5] <= img[6395];\
        in_img_array[14][21][6] <= img[6396];\
        in_img_array[14][21][7] <= img[6397];\
        in_img_array[14][21][8] <= img[6398];\
        in_img_array[14][21][9] <= img[6399];\
        in_img_array[14][21][10] <= img[6400];\
        in_img_array[14][21][11] <= img[6401];\
        in_img_array[14][21][12] <= img[6402];\
        in_img_array[14][21][13] <= img[6403];\
        in_img_array[14][21][14] <= img[6404];\
        in_img_array[14][21][15] <= img[6405];\
        in_img_array[14][21][16] <= img[6406];\
        in_img_array[14][21][17] <= img[6407];\
        in_img_array[14][22][0] <= img[6408];\
        in_img_array[14][22][1] <= img[6409];\
        in_img_array[14][22][2] <= img[6410];\
        in_img_array[14][22][3] <= img[6411];\
        in_img_array[14][22][4] <= img[6412];\
        in_img_array[14][22][5] <= img[6413];\
        in_img_array[14][22][6] <= img[6414];\
        in_img_array[14][22][7] <= img[6415];\
        in_img_array[14][22][8] <= img[6416];\
        in_img_array[14][22][9] <= img[6417];\
        in_img_array[14][22][10] <= img[6418];\
        in_img_array[14][22][11] <= img[6419];\
        in_img_array[14][22][12] <= img[6420];\
        in_img_array[14][22][13] <= img[6421];\
        in_img_array[14][22][14] <= img[6422];\
        in_img_array[14][22][15] <= img[6423];\
        in_img_array[14][22][16] <= img[6424];\
        in_img_array[14][22][17] <= img[6425];\
        in_img_array[14][23][0] <= img[6426];\
        in_img_array[14][23][1] <= img[6427];\
        in_img_array[14][23][2] <= img[6428];\
        in_img_array[14][23][3] <= img[6429];\
        in_img_array[14][23][4] <= img[6430];\
        in_img_array[14][23][5] <= img[6431];\
        in_img_array[14][23][6] <= img[6432];\
        in_img_array[14][23][7] <= img[6433];\
        in_img_array[14][23][8] <= img[6434];\
        in_img_array[14][23][9] <= img[6435];\
        in_img_array[14][23][10] <= img[6436];\
        in_img_array[14][23][11] <= img[6437];\
        in_img_array[14][23][12] <= img[6438];\
        in_img_array[14][23][13] <= img[6439];\
        in_img_array[14][23][14] <= img[6440];\
        in_img_array[14][23][15] <= img[6441];\
        in_img_array[14][23][16] <= img[6442];\
        in_img_array[14][23][17] <= img[6443];\
        in_img_array[14][24][0] <= img[6444];\
        in_img_array[14][24][1] <= img[6445];\
        in_img_array[14][24][2] <= img[6446];\
        in_img_array[14][24][3] <= img[6447];\
        in_img_array[14][24][4] <= img[6448];\
        in_img_array[14][24][5] <= img[6449];\
        in_img_array[14][24][6] <= img[6450];\
        in_img_array[14][24][7] <= img[6451];\
        in_img_array[14][24][8] <= img[6452];\
        in_img_array[14][24][9] <= img[6453];\
        in_img_array[14][24][10] <= img[6454];\
        in_img_array[14][24][11] <= img[6455];\
        in_img_array[14][24][12] <= img[6456];\
        in_img_array[14][24][13] <= img[6457];\
        in_img_array[14][24][14] <= img[6458];\
        in_img_array[14][24][15] <= img[6459];\
        in_img_array[14][24][16] <= img[6460];\
        in_img_array[14][24][17] <= img[6461];\
        in_img_array[14][25][0] <= img[6462];\
        in_img_array[14][25][1] <= img[6463];\
        in_img_array[14][25][2] <= img[6464];\
        in_img_array[14][25][3] <= img[6465];\
        in_img_array[14][25][4] <= img[6466];\
        in_img_array[14][25][5] <= img[6467];\
        in_img_array[14][25][6] <= img[6468];\
        in_img_array[14][25][7] <= img[6469];\
        in_img_array[14][25][8] <= img[6470];\
        in_img_array[14][25][9] <= img[6471];\
        in_img_array[14][25][10] <= img[6472];\
        in_img_array[14][25][11] <= img[6473];\
        in_img_array[14][25][12] <= img[6474];\
        in_img_array[14][25][13] <= img[6475];\
        in_img_array[14][25][14] <= img[6476];\
        in_img_array[14][25][15] <= img[6477];\
        in_img_array[14][25][16] <= img[6478];\
        in_img_array[14][25][17] <= img[6479];\
        in_img_array[14][26][0] <= img[6480];\
        in_img_array[14][26][1] <= img[6481];\
        in_img_array[14][26][2] <= img[6482];\
        in_img_array[14][26][3] <= img[6483];\
        in_img_array[14][26][4] <= img[6484];\
        in_img_array[14][26][5] <= img[6485];\
        in_img_array[14][26][6] <= img[6486];\
        in_img_array[14][26][7] <= img[6487];\
        in_img_array[14][26][8] <= img[6488];\
        in_img_array[14][26][9] <= img[6489];\
        in_img_array[14][26][10] <= img[6490];\
        in_img_array[14][26][11] <= img[6491];\
        in_img_array[14][26][12] <= img[6492];\
        in_img_array[14][26][13] <= img[6493];\
        in_img_array[14][26][14] <= img[6494];\
        in_img_array[14][26][15] <= img[6495];\
        in_img_array[14][26][16] <= img[6496];\
        in_img_array[14][26][17] <= img[6497];\
        in_img_array[14][27][0] <= img[6498];\
        in_img_array[14][27][1] <= img[6499];\
        in_img_array[14][27][2] <= img[6500];\
        in_img_array[14][27][3] <= img[6501];\
        in_img_array[14][27][4] <= img[6502];\
        in_img_array[14][27][5] <= img[6503];\
        in_img_array[14][27][6] <= img[6504];\
        in_img_array[14][27][7] <= img[6505];\
        in_img_array[14][27][8] <= img[6506];\
        in_img_array[14][27][9] <= img[6507];\
        in_img_array[14][27][10] <= img[6508];\
        in_img_array[14][27][11] <= img[6509];\
        in_img_array[14][27][12] <= img[6510];\
        in_img_array[14][27][13] <= img[6511];\
        in_img_array[14][27][14] <= img[6512];\
        in_img_array[14][27][15] <= img[6513];\
        in_img_array[14][27][16] <= img[6514];\
        in_img_array[14][27][17] <= img[6515];\
        in_img_array[14][28][0] <= img[6516];\
        in_img_array[14][28][1] <= img[6517];\
        in_img_array[14][28][2] <= img[6518];\
        in_img_array[14][28][3] <= img[6519];\
        in_img_array[14][28][4] <= img[6520];\
        in_img_array[14][28][5] <= img[6521];\
        in_img_array[14][28][6] <= img[6522];\
        in_img_array[14][28][7] <= img[6523];\
        in_img_array[14][28][8] <= img[6524];\
        in_img_array[14][28][9] <= img[6525];\
        in_img_array[14][28][10] <= img[6526];\
        in_img_array[14][28][11] <= img[6527];\
        in_img_array[14][28][12] <= img[6528];\
        in_img_array[14][28][13] <= img[6529];\
        in_img_array[14][28][14] <= img[6530];\
        in_img_array[14][28][15] <= img[6531];\
        in_img_array[14][28][16] <= img[6532];\
        in_img_array[14][28][17] <= img[6533];\
        in_img_array[14][29][0] <= img[6534];\
        in_img_array[14][29][1] <= img[6535];\
        in_img_array[14][29][2] <= img[6536];\
        in_img_array[14][29][3] <= img[6537];\
        in_img_array[14][29][4] <= img[6538];\
        in_img_array[14][29][5] <= img[6539];\
        in_img_array[14][29][6] <= img[6540];\
        in_img_array[14][29][7] <= img[6541];\
        in_img_array[14][29][8] <= img[6542];\
        in_img_array[14][29][9] <= img[6543];\
        in_img_array[14][29][10] <= img[6544];\
        in_img_array[14][29][11] <= img[6545];\
        in_img_array[14][29][12] <= img[6546];\
        in_img_array[14][29][13] <= img[6547];\
        in_img_array[14][29][14] <= img[6548];\
        in_img_array[14][29][15] <= img[6549];\
        in_img_array[14][29][16] <= img[6550];\
        in_img_array[14][29][17] <= img[6551];\
        in_img_array[15][2][0] <= img[6552];\
        in_img_array[15][2][1] <= img[6553];\
        in_img_array[15][2][2] <= img[6554];\
        in_img_array[15][2][3] <= img[6555];\
        in_img_array[15][2][4] <= img[6556];\
        in_img_array[15][2][5] <= img[6557];\
        in_img_array[15][2][6] <= img[6558];\
        in_img_array[15][2][7] <= img[6559];\
        in_img_array[15][2][8] <= img[6560];\
        in_img_array[15][2][9] <= img[6561];\
        in_img_array[15][2][10] <= img[6562];\
        in_img_array[15][2][11] <= img[6563];\
        in_img_array[15][2][12] <= img[6564];\
        in_img_array[15][2][13] <= img[6565];\
        in_img_array[15][2][14] <= img[6566];\
        in_img_array[15][2][15] <= img[6567];\
        in_img_array[15][2][16] <= img[6568];\
        in_img_array[15][2][17] <= img[6569];\
        in_img_array[15][3][0] <= img[6570];\
        in_img_array[15][3][1] <= img[6571];\
        in_img_array[15][3][2] <= img[6572];\
        in_img_array[15][3][3] <= img[6573];\
        in_img_array[15][3][4] <= img[6574];\
        in_img_array[15][3][5] <= img[6575];\
        in_img_array[15][3][6] <= img[6576];\
        in_img_array[15][3][7] <= img[6577];\
        in_img_array[15][3][8] <= img[6578];\
        in_img_array[15][3][9] <= img[6579];\
        in_img_array[15][3][10] <= img[6580];\
        in_img_array[15][3][11] <= img[6581];\
        in_img_array[15][3][12] <= img[6582];\
        in_img_array[15][3][13] <= img[6583];\
        in_img_array[15][3][14] <= img[6584];\
        in_img_array[15][3][15] <= img[6585];\
        in_img_array[15][3][16] <= img[6586];\
        in_img_array[15][3][17] <= img[6587];\
        in_img_array[15][4][0] <= img[6588];\
        in_img_array[15][4][1] <= img[6589];\
        in_img_array[15][4][2] <= img[6590];\
        in_img_array[15][4][3] <= img[6591];\
        in_img_array[15][4][4] <= img[6592];\
        in_img_array[15][4][5] <= img[6593];\
        in_img_array[15][4][6] <= img[6594];\
        in_img_array[15][4][7] <= img[6595];\
        in_img_array[15][4][8] <= img[6596];\
        in_img_array[15][4][9] <= img[6597];\
        in_img_array[15][4][10] <= img[6598];\
        in_img_array[15][4][11] <= img[6599];\
        in_img_array[15][4][12] <= img[6600];\
        in_img_array[15][4][13] <= img[6601];\
        in_img_array[15][4][14] <= img[6602];\
        in_img_array[15][4][15] <= img[6603];\
        in_img_array[15][4][16] <= img[6604];\
        in_img_array[15][4][17] <= img[6605];\
        in_img_array[15][5][0] <= img[6606];\
        in_img_array[15][5][1] <= img[6607];\
        in_img_array[15][5][2] <= img[6608];\
        in_img_array[15][5][3] <= img[6609];\
        in_img_array[15][5][4] <= img[6610];\
        in_img_array[15][5][5] <= img[6611];\
        in_img_array[15][5][6] <= img[6612];\
        in_img_array[15][5][7] <= img[6613];\
        in_img_array[15][5][8] <= img[6614];\
        in_img_array[15][5][9] <= img[6615];\
        in_img_array[15][5][10] <= img[6616];\
        in_img_array[15][5][11] <= img[6617];\
        in_img_array[15][5][12] <= img[6618];\
        in_img_array[15][5][13] <= img[6619];\
        in_img_array[15][5][14] <= img[6620];\
        in_img_array[15][5][15] <= img[6621];\
        in_img_array[15][5][16] <= img[6622];\
        in_img_array[15][5][17] <= img[6623];\
        in_img_array[15][6][0] <= img[6624];\
        in_img_array[15][6][1] <= img[6625];\
        in_img_array[15][6][2] <= img[6626];\
        in_img_array[15][6][3] <= img[6627];\
        in_img_array[15][6][4] <= img[6628];\
        in_img_array[15][6][5] <= img[6629];\
        in_img_array[15][6][6] <= img[6630];\
        in_img_array[15][6][7] <= img[6631];\
        in_img_array[15][6][8] <= img[6632];\
        in_img_array[15][6][9] <= img[6633];\
        in_img_array[15][6][10] <= img[6634];\
        in_img_array[15][6][11] <= img[6635];\
        in_img_array[15][6][12] <= img[6636];\
        in_img_array[15][6][13] <= img[6637];\
        in_img_array[15][6][14] <= img[6638];\
        in_img_array[15][6][15] <= img[6639];\
        in_img_array[15][6][16] <= img[6640];\
        in_img_array[15][6][17] <= img[6641];\
        in_img_array[15][7][0] <= img[6642];\
        in_img_array[15][7][1] <= img[6643];\
        in_img_array[15][7][2] <= img[6644];\
        in_img_array[15][7][3] <= img[6645];\
        in_img_array[15][7][4] <= img[6646];\
        in_img_array[15][7][5] <= img[6647];\
        in_img_array[15][7][6] <= img[6648];\
        in_img_array[15][7][7] <= img[6649];\
        in_img_array[15][7][8] <= img[6650];\
        in_img_array[15][7][9] <= img[6651];\
        in_img_array[15][7][10] <= img[6652];\
        in_img_array[15][7][11] <= img[6653];\
        in_img_array[15][7][12] <= img[6654];\
        in_img_array[15][7][13] <= img[6655];\
        in_img_array[15][7][14] <= img[6656];\
        in_img_array[15][7][15] <= img[6657];\
        in_img_array[15][7][16] <= img[6658];\
        in_img_array[15][7][17] <= img[6659];\
        in_img_array[15][8][0] <= img[6660];\
        in_img_array[15][8][1] <= img[6661];\
        in_img_array[15][8][2] <= img[6662];\
        in_img_array[15][8][3] <= img[6663];\
        in_img_array[15][8][4] <= img[6664];\
        in_img_array[15][8][5] <= img[6665];\
        in_img_array[15][8][6] <= img[6666];\
        in_img_array[15][8][7] <= img[6667];\
        in_img_array[15][8][8] <= img[6668];\
        in_img_array[15][8][9] <= img[6669];\
        in_img_array[15][8][10] <= img[6670];\
        in_img_array[15][8][11] <= img[6671];\
        in_img_array[15][8][12] <= img[6672];\
        in_img_array[15][8][13] <= img[6673];\
        in_img_array[15][8][14] <= img[6674];\
        in_img_array[15][8][15] <= img[6675];\
        in_img_array[15][8][16] <= img[6676];\
        in_img_array[15][8][17] <= img[6677];\
        in_img_array[15][9][0] <= img[6678];\
        in_img_array[15][9][1] <= img[6679];\
        in_img_array[15][9][2] <= img[6680];\
        in_img_array[15][9][3] <= img[6681];\
        in_img_array[15][9][4] <= img[6682];\
        in_img_array[15][9][5] <= img[6683];\
        in_img_array[15][9][6] <= img[6684];\
        in_img_array[15][9][7] <= img[6685];\
        in_img_array[15][9][8] <= img[6686];\
        in_img_array[15][9][9] <= img[6687];\
        in_img_array[15][9][10] <= img[6688];\
        in_img_array[15][9][11] <= img[6689];\
        in_img_array[15][9][12] <= img[6690];\
        in_img_array[15][9][13] <= img[6691];\
        in_img_array[15][9][14] <= img[6692];\
        in_img_array[15][9][15] <= img[6693];\
        in_img_array[15][9][16] <= img[6694];\
        in_img_array[15][9][17] <= img[6695];\
        in_img_array[15][10][0] <= img[6696];\
        in_img_array[15][10][1] <= img[6697];\
        in_img_array[15][10][2] <= img[6698];\
        in_img_array[15][10][3] <= img[6699];\
        in_img_array[15][10][4] <= img[6700];\
        in_img_array[15][10][5] <= img[6701];\
        in_img_array[15][10][6] <= img[6702];\
        in_img_array[15][10][7] <= img[6703];\
        in_img_array[15][10][8] <= img[6704];\
        in_img_array[15][10][9] <= img[6705];\
        in_img_array[15][10][10] <= img[6706];\
        in_img_array[15][10][11] <= img[6707];\
        in_img_array[15][10][12] <= img[6708];\
        in_img_array[15][10][13] <= img[6709];\
        in_img_array[15][10][14] <= img[6710];\
        in_img_array[15][10][15] <= img[6711];\
        in_img_array[15][10][16] <= img[6712];\
        in_img_array[15][10][17] <= img[6713];\
        in_img_array[15][11][0] <= img[6714];\
        in_img_array[15][11][1] <= img[6715];\
        in_img_array[15][11][2] <= img[6716];\
        in_img_array[15][11][3] <= img[6717];\
        in_img_array[15][11][4] <= img[6718];\
        in_img_array[15][11][5] <= img[6719];\
        in_img_array[15][11][6] <= img[6720];\
        in_img_array[15][11][7] <= img[6721];\
        in_img_array[15][11][8] <= img[6722];\
        in_img_array[15][11][9] <= img[6723];\
        in_img_array[15][11][10] <= img[6724];\
        in_img_array[15][11][11] <= img[6725];\
        in_img_array[15][11][12] <= img[6726];\
        in_img_array[15][11][13] <= img[6727];\
        in_img_array[15][11][14] <= img[6728];\
        in_img_array[15][11][15] <= img[6729];\
        in_img_array[15][11][16] <= img[6730];\
        in_img_array[15][11][17] <= img[6731];\
        in_img_array[15][12][0] <= img[6732];\
        in_img_array[15][12][1] <= img[6733];\
        in_img_array[15][12][2] <= img[6734];\
        in_img_array[15][12][3] <= img[6735];\
        in_img_array[15][12][4] <= img[6736];\
        in_img_array[15][12][5] <= img[6737];\
        in_img_array[15][12][6] <= img[6738];\
        in_img_array[15][12][7] <= img[6739];\
        in_img_array[15][12][8] <= img[6740];\
        in_img_array[15][12][9] <= img[6741];\
        in_img_array[15][12][10] <= img[6742];\
        in_img_array[15][12][11] <= img[6743];\
        in_img_array[15][12][12] <= img[6744];\
        in_img_array[15][12][13] <= img[6745];\
        in_img_array[15][12][14] <= img[6746];\
        in_img_array[15][12][15] <= img[6747];\
        in_img_array[15][12][16] <= img[6748];\
        in_img_array[15][12][17] <= img[6749];\
        in_img_array[15][13][0] <= img[6750];\
        in_img_array[15][13][1] <= img[6751];\
        in_img_array[15][13][2] <= img[6752];\
        in_img_array[15][13][3] <= img[6753];\
        in_img_array[15][13][4] <= img[6754];\
        in_img_array[15][13][5] <= img[6755];\
        in_img_array[15][13][6] <= img[6756];\
        in_img_array[15][13][7] <= img[6757];\
        in_img_array[15][13][8] <= img[6758];\
        in_img_array[15][13][9] <= img[6759];\
        in_img_array[15][13][10] <= img[6760];\
        in_img_array[15][13][11] <= img[6761];\
        in_img_array[15][13][12] <= img[6762];\
        in_img_array[15][13][13] <= img[6763];\
        in_img_array[15][13][14] <= img[6764];\
        in_img_array[15][13][15] <= img[6765];\
        in_img_array[15][13][16] <= img[6766];\
        in_img_array[15][13][17] <= img[6767];\
        in_img_array[15][14][0] <= img[6768];\
        in_img_array[15][14][1] <= img[6769];\
        in_img_array[15][14][2] <= img[6770];\
        in_img_array[15][14][3] <= img[6771];\
        in_img_array[15][14][4] <= img[6772];\
        in_img_array[15][14][5] <= img[6773];\
        in_img_array[15][14][6] <= img[6774];\
        in_img_array[15][14][7] <= img[6775];\
        in_img_array[15][14][8] <= img[6776];\
        in_img_array[15][14][9] <= img[6777];\
        in_img_array[15][14][10] <= img[6778];\
        in_img_array[15][14][11] <= img[6779];\
        in_img_array[15][14][12] <= img[6780];\
        in_img_array[15][14][13] <= img[6781];\
        in_img_array[15][14][14] <= img[6782];\
        in_img_array[15][14][15] <= img[6783];\
        in_img_array[15][14][16] <= img[6784];\
        in_img_array[15][14][17] <= img[6785];\
        in_img_array[15][15][0] <= img[6786];\
        in_img_array[15][15][1] <= img[6787];\
        in_img_array[15][15][2] <= img[6788];\
        in_img_array[15][15][3] <= img[6789];\
        in_img_array[15][15][4] <= img[6790];\
        in_img_array[15][15][5] <= img[6791];\
        in_img_array[15][15][6] <= img[6792];\
        in_img_array[15][15][7] <= img[6793];\
        in_img_array[15][15][8] <= img[6794];\
        in_img_array[15][15][9] <= img[6795];\
        in_img_array[15][15][10] <= img[6796];\
        in_img_array[15][15][11] <= img[6797];\
        in_img_array[15][15][12] <= img[6798];\
        in_img_array[15][15][13] <= img[6799];\
        in_img_array[15][15][14] <= img[6800];\
        in_img_array[15][15][15] <= img[6801];\
        in_img_array[15][15][16] <= img[6802];\
        in_img_array[15][15][17] <= img[6803];\
        in_img_array[15][16][0] <= img[6804];\
        in_img_array[15][16][1] <= img[6805];\
        in_img_array[15][16][2] <= img[6806];\
        in_img_array[15][16][3] <= img[6807];\
        in_img_array[15][16][4] <= img[6808];\
        in_img_array[15][16][5] <= img[6809];\
        in_img_array[15][16][6] <= img[6810];\
        in_img_array[15][16][7] <= img[6811];\
        in_img_array[15][16][8] <= img[6812];\
        in_img_array[15][16][9] <= img[6813];\
        in_img_array[15][16][10] <= img[6814];\
        in_img_array[15][16][11] <= img[6815];\
        in_img_array[15][16][12] <= img[6816];\
        in_img_array[15][16][13] <= img[6817];\
        in_img_array[15][16][14] <= img[6818];\
        in_img_array[15][16][15] <= img[6819];\
        in_img_array[15][16][16] <= img[6820];\
        in_img_array[15][16][17] <= img[6821];\
        in_img_array[15][17][0] <= img[6822];\
        in_img_array[15][17][1] <= img[6823];\
        in_img_array[15][17][2] <= img[6824];\
        in_img_array[15][17][3] <= img[6825];\
        in_img_array[15][17][4] <= img[6826];\
        in_img_array[15][17][5] <= img[6827];\
        in_img_array[15][17][6] <= img[6828];\
        in_img_array[15][17][7] <= img[6829];\
        in_img_array[15][17][8] <= img[6830];\
        in_img_array[15][17][9] <= img[6831];\
        in_img_array[15][17][10] <= img[6832];\
        in_img_array[15][17][11] <= img[6833];\
        in_img_array[15][17][12] <= img[6834];\
        in_img_array[15][17][13] <= img[6835];\
        in_img_array[15][17][14] <= img[6836];\
        in_img_array[15][17][15] <= img[6837];\
        in_img_array[15][17][16] <= img[6838];\
        in_img_array[15][17][17] <= img[6839];\
        in_img_array[15][18][0] <= img[6840];\
        in_img_array[15][18][1] <= img[6841];\
        in_img_array[15][18][2] <= img[6842];\
        in_img_array[15][18][3] <= img[6843];\
        in_img_array[15][18][4] <= img[6844];\
        in_img_array[15][18][5] <= img[6845];\
        in_img_array[15][18][6] <= img[6846];\
        in_img_array[15][18][7] <= img[6847];\
        in_img_array[15][18][8] <= img[6848];\
        in_img_array[15][18][9] <= img[6849];\
        in_img_array[15][18][10] <= img[6850];\
        in_img_array[15][18][11] <= img[6851];\
        in_img_array[15][18][12] <= img[6852];\
        in_img_array[15][18][13] <= img[6853];\
        in_img_array[15][18][14] <= img[6854];\
        in_img_array[15][18][15] <= img[6855];\
        in_img_array[15][18][16] <= img[6856];\
        in_img_array[15][18][17] <= img[6857];\
        in_img_array[15][19][0] <= img[6858];\
        in_img_array[15][19][1] <= img[6859];\
        in_img_array[15][19][2] <= img[6860];\
        in_img_array[15][19][3] <= img[6861];\
        in_img_array[15][19][4] <= img[6862];\
        in_img_array[15][19][5] <= img[6863];\
        in_img_array[15][19][6] <= img[6864];\
        in_img_array[15][19][7] <= img[6865];\
        in_img_array[15][19][8] <= img[6866];\
        in_img_array[15][19][9] <= img[6867];\
        in_img_array[15][19][10] <= img[6868];\
        in_img_array[15][19][11] <= img[6869];\
        in_img_array[15][19][12] <= img[6870];\
        in_img_array[15][19][13] <= img[6871];\
        in_img_array[15][19][14] <= img[6872];\
        in_img_array[15][19][15] <= img[6873];\
        in_img_array[15][19][16] <= img[6874];\
        in_img_array[15][19][17] <= img[6875];\
        in_img_array[15][20][0] <= img[6876];\
        in_img_array[15][20][1] <= img[6877];\
        in_img_array[15][20][2] <= img[6878];\
        in_img_array[15][20][3] <= img[6879];\
        in_img_array[15][20][4] <= img[6880];\
        in_img_array[15][20][5] <= img[6881];\
        in_img_array[15][20][6] <= img[6882];\
        in_img_array[15][20][7] <= img[6883];\
        in_img_array[15][20][8] <= img[6884];\
        in_img_array[15][20][9] <= img[6885];\
        in_img_array[15][20][10] <= img[6886];\
        in_img_array[15][20][11] <= img[6887];\
        in_img_array[15][20][12] <= img[6888];\
        in_img_array[15][20][13] <= img[6889];\
        in_img_array[15][20][14] <= img[6890];\
        in_img_array[15][20][15] <= img[6891];\
        in_img_array[15][20][16] <= img[6892];\
        in_img_array[15][20][17] <= img[6893];\
        in_img_array[15][21][0] <= img[6894];\
        in_img_array[15][21][1] <= img[6895];\
        in_img_array[15][21][2] <= img[6896];\
        in_img_array[15][21][3] <= img[6897];\
        in_img_array[15][21][4] <= img[6898];\
        in_img_array[15][21][5] <= img[6899];\
        in_img_array[15][21][6] <= img[6900];\
        in_img_array[15][21][7] <= img[6901];\
        in_img_array[15][21][8] <= img[6902];\
        in_img_array[15][21][9] <= img[6903];\
        in_img_array[15][21][10] <= img[6904];\
        in_img_array[15][21][11] <= img[6905];\
        in_img_array[15][21][12] <= img[6906];\
        in_img_array[15][21][13] <= img[6907];\
        in_img_array[15][21][14] <= img[6908];\
        in_img_array[15][21][15] <= img[6909];\
        in_img_array[15][21][16] <= img[6910];\
        in_img_array[15][21][17] <= img[6911];\
        in_img_array[15][22][0] <= img[6912];\
        in_img_array[15][22][1] <= img[6913];\
        in_img_array[15][22][2] <= img[6914];\
        in_img_array[15][22][3] <= img[6915];\
        in_img_array[15][22][4] <= img[6916];\
        in_img_array[15][22][5] <= img[6917];\
        in_img_array[15][22][6] <= img[6918];\
        in_img_array[15][22][7] <= img[6919];\
        in_img_array[15][22][8] <= img[6920];\
        in_img_array[15][22][9] <= img[6921];\
        in_img_array[15][22][10] <= img[6922];\
        in_img_array[15][22][11] <= img[6923];\
        in_img_array[15][22][12] <= img[6924];\
        in_img_array[15][22][13] <= img[6925];\
        in_img_array[15][22][14] <= img[6926];\
        in_img_array[15][22][15] <= img[6927];\
        in_img_array[15][22][16] <= img[6928];\
        in_img_array[15][22][17] <= img[6929];\
        in_img_array[15][23][0] <= img[6930];\
        in_img_array[15][23][1] <= img[6931];\
        in_img_array[15][23][2] <= img[6932];\
        in_img_array[15][23][3] <= img[6933];\
        in_img_array[15][23][4] <= img[6934];\
        in_img_array[15][23][5] <= img[6935];\
        in_img_array[15][23][6] <= img[6936];\
        in_img_array[15][23][7] <= img[6937];\
        in_img_array[15][23][8] <= img[6938];\
        in_img_array[15][23][9] <= img[6939];\
        in_img_array[15][23][10] <= img[6940];\
        in_img_array[15][23][11] <= img[6941];\
        in_img_array[15][23][12] <= img[6942];\
        in_img_array[15][23][13] <= img[6943];\
        in_img_array[15][23][14] <= img[6944];\
        in_img_array[15][23][15] <= img[6945];\
        in_img_array[15][23][16] <= img[6946];\
        in_img_array[15][23][17] <= img[6947];\
        in_img_array[15][24][0] <= img[6948];\
        in_img_array[15][24][1] <= img[6949];\
        in_img_array[15][24][2] <= img[6950];\
        in_img_array[15][24][3] <= img[6951];\
        in_img_array[15][24][4] <= img[6952];\
        in_img_array[15][24][5] <= img[6953];\
        in_img_array[15][24][6] <= img[6954];\
        in_img_array[15][24][7] <= img[6955];\
        in_img_array[15][24][8] <= img[6956];\
        in_img_array[15][24][9] <= img[6957];\
        in_img_array[15][24][10] <= img[6958];\
        in_img_array[15][24][11] <= img[6959];\
        in_img_array[15][24][12] <= img[6960];\
        in_img_array[15][24][13] <= img[6961];\
        in_img_array[15][24][14] <= img[6962];\
        in_img_array[15][24][15] <= img[6963];\
        in_img_array[15][24][16] <= img[6964];\
        in_img_array[15][24][17] <= img[6965];\
        in_img_array[15][25][0] <= img[6966];\
        in_img_array[15][25][1] <= img[6967];\
        in_img_array[15][25][2] <= img[6968];\
        in_img_array[15][25][3] <= img[6969];\
        in_img_array[15][25][4] <= img[6970];\
        in_img_array[15][25][5] <= img[6971];\
        in_img_array[15][25][6] <= img[6972];\
        in_img_array[15][25][7] <= img[6973];\
        in_img_array[15][25][8] <= img[6974];\
        in_img_array[15][25][9] <= img[6975];\
        in_img_array[15][25][10] <= img[6976];\
        in_img_array[15][25][11] <= img[6977];\
        in_img_array[15][25][12] <= img[6978];\
        in_img_array[15][25][13] <= img[6979];\
        in_img_array[15][25][14] <= img[6980];\
        in_img_array[15][25][15] <= img[6981];\
        in_img_array[15][25][16] <= img[6982];\
        in_img_array[15][25][17] <= img[6983];\
        in_img_array[15][26][0] <= img[6984];\
        in_img_array[15][26][1] <= img[6985];\
        in_img_array[15][26][2] <= img[6986];\
        in_img_array[15][26][3] <= img[6987];\
        in_img_array[15][26][4] <= img[6988];\
        in_img_array[15][26][5] <= img[6989];\
        in_img_array[15][26][6] <= img[6990];\
        in_img_array[15][26][7] <= img[6991];\
        in_img_array[15][26][8] <= img[6992];\
        in_img_array[15][26][9] <= img[6993];\
        in_img_array[15][26][10] <= img[6994];\
        in_img_array[15][26][11] <= img[6995];\
        in_img_array[15][26][12] <= img[6996];\
        in_img_array[15][26][13] <= img[6997];\
        in_img_array[15][26][14] <= img[6998];\
        in_img_array[15][26][15] <= img[6999];\
        in_img_array[15][26][16] <= img[7000];\
        in_img_array[15][26][17] <= img[7001];\
        in_img_array[15][27][0] <= img[7002];\
        in_img_array[15][27][1] <= img[7003];\
        in_img_array[15][27][2] <= img[7004];\
        in_img_array[15][27][3] <= img[7005];\
        in_img_array[15][27][4] <= img[7006];\
        in_img_array[15][27][5] <= img[7007];\
        in_img_array[15][27][6] <= img[7008];\
        in_img_array[15][27][7] <= img[7009];\
        in_img_array[15][27][8] <= img[7010];\
        in_img_array[15][27][9] <= img[7011];\
        in_img_array[15][27][10] <= img[7012];\
        in_img_array[15][27][11] <= img[7013];\
        in_img_array[15][27][12] <= img[7014];\
        in_img_array[15][27][13] <= img[7015];\
        in_img_array[15][27][14] <= img[7016];\
        in_img_array[15][27][15] <= img[7017];\
        in_img_array[15][27][16] <= img[7018];\
        in_img_array[15][27][17] <= img[7019];\
        in_img_array[15][28][0] <= img[7020];\
        in_img_array[15][28][1] <= img[7021];\
        in_img_array[15][28][2] <= img[7022];\
        in_img_array[15][28][3] <= img[7023];\
        in_img_array[15][28][4] <= img[7024];\
        in_img_array[15][28][5] <= img[7025];\
        in_img_array[15][28][6] <= img[7026];\
        in_img_array[15][28][7] <= img[7027];\
        in_img_array[15][28][8] <= img[7028];\
        in_img_array[15][28][9] <= img[7029];\
        in_img_array[15][28][10] <= img[7030];\
        in_img_array[15][28][11] <= img[7031];\
        in_img_array[15][28][12] <= img[7032];\
        in_img_array[15][28][13] <= img[7033];\
        in_img_array[15][28][14] <= img[7034];\
        in_img_array[15][28][15] <= img[7035];\
        in_img_array[15][28][16] <= img[7036];\
        in_img_array[15][28][17] <= img[7037];\
        in_img_array[15][29][0] <= img[7038];\
        in_img_array[15][29][1] <= img[7039];\
        in_img_array[15][29][2] <= img[7040];\
        in_img_array[15][29][3] <= img[7041];\
        in_img_array[15][29][4] <= img[7042];\
        in_img_array[15][29][5] <= img[7043];\
        in_img_array[15][29][6] <= img[7044];\
        in_img_array[15][29][7] <= img[7045];\
        in_img_array[15][29][8] <= img[7046];\
        in_img_array[15][29][9] <= img[7047];\
        in_img_array[15][29][10] <= img[7048];\
        in_img_array[15][29][11] <= img[7049];\
        in_img_array[15][29][12] <= img[7050];\
        in_img_array[15][29][13] <= img[7051];\
        in_img_array[15][29][14] <= img[7052];\
        in_img_array[15][29][15] <= img[7053];\
        in_img_array[15][29][16] <= img[7054];\
        in_img_array[15][29][17] <= img[7055];\
        in_img_array[16][2][0] <= img[7056];\
        in_img_array[16][2][1] <= img[7057];\
        in_img_array[16][2][2] <= img[7058];\
        in_img_array[16][2][3] <= img[7059];\
        in_img_array[16][2][4] <= img[7060];\
        in_img_array[16][2][5] <= img[7061];\
        in_img_array[16][2][6] <= img[7062];\
        in_img_array[16][2][7] <= img[7063];\
        in_img_array[16][2][8] <= img[7064];\
        in_img_array[16][2][9] <= img[7065];\
        in_img_array[16][2][10] <= img[7066];\
        in_img_array[16][2][11] <= img[7067];\
        in_img_array[16][2][12] <= img[7068];\
        in_img_array[16][2][13] <= img[7069];\
        in_img_array[16][2][14] <= img[7070];\
        in_img_array[16][2][15] <= img[7071];\
        in_img_array[16][2][16] <= img[7072];\
        in_img_array[16][2][17] <= img[7073];\
        in_img_array[16][3][0] <= img[7074];\
        in_img_array[16][3][1] <= img[7075];\
        in_img_array[16][3][2] <= img[7076];\
        in_img_array[16][3][3] <= img[7077];\
        in_img_array[16][3][4] <= img[7078];\
        in_img_array[16][3][5] <= img[7079];\
        in_img_array[16][3][6] <= img[7080];\
        in_img_array[16][3][7] <= img[7081];\
        in_img_array[16][3][8] <= img[7082];\
        in_img_array[16][3][9] <= img[7083];\
        in_img_array[16][3][10] <= img[7084];\
        in_img_array[16][3][11] <= img[7085];\
        in_img_array[16][3][12] <= img[7086];\
        in_img_array[16][3][13] <= img[7087];\
        in_img_array[16][3][14] <= img[7088];\
        in_img_array[16][3][15] <= img[7089];\
        in_img_array[16][3][16] <= img[7090];\
        in_img_array[16][3][17] <= img[7091];\
        in_img_array[16][4][0] <= img[7092];\
        in_img_array[16][4][1] <= img[7093];\
        in_img_array[16][4][2] <= img[7094];\
        in_img_array[16][4][3] <= img[7095];\
        in_img_array[16][4][4] <= img[7096];\
        in_img_array[16][4][5] <= img[7097];\
        in_img_array[16][4][6] <= img[7098];\
        in_img_array[16][4][7] <= img[7099];\
        in_img_array[16][4][8] <= img[7100];\
        in_img_array[16][4][9] <= img[7101];\
        in_img_array[16][4][10] <= img[7102];\
        in_img_array[16][4][11] <= img[7103];\
        in_img_array[16][4][12] <= img[7104];\
        in_img_array[16][4][13] <= img[7105];\
        in_img_array[16][4][14] <= img[7106];\
        in_img_array[16][4][15] <= img[7107];\
        in_img_array[16][4][16] <= img[7108];\
        in_img_array[16][4][17] <= img[7109];\
        in_img_array[16][5][0] <= img[7110];\
        in_img_array[16][5][1] <= img[7111];\
        in_img_array[16][5][2] <= img[7112];\
        in_img_array[16][5][3] <= img[7113];\
        in_img_array[16][5][4] <= img[7114];\
        in_img_array[16][5][5] <= img[7115];\
        in_img_array[16][5][6] <= img[7116];\
        in_img_array[16][5][7] <= img[7117];\
        in_img_array[16][5][8] <= img[7118];\
        in_img_array[16][5][9] <= img[7119];\
        in_img_array[16][5][10] <= img[7120];\
        in_img_array[16][5][11] <= img[7121];\
        in_img_array[16][5][12] <= img[7122];\
        in_img_array[16][5][13] <= img[7123];\
        in_img_array[16][5][14] <= img[7124];\
        in_img_array[16][5][15] <= img[7125];\
        in_img_array[16][5][16] <= img[7126];\
        in_img_array[16][5][17] <= img[7127];\
        in_img_array[16][6][0] <= img[7128];\
        in_img_array[16][6][1] <= img[7129];\
        in_img_array[16][6][2] <= img[7130];\
        in_img_array[16][6][3] <= img[7131];\
        in_img_array[16][6][4] <= img[7132];\
        in_img_array[16][6][5] <= img[7133];\
        in_img_array[16][6][6] <= img[7134];\
        in_img_array[16][6][7] <= img[7135];\
        in_img_array[16][6][8] <= img[7136];\
        in_img_array[16][6][9] <= img[7137];\
        in_img_array[16][6][10] <= img[7138];\
        in_img_array[16][6][11] <= img[7139];\
        in_img_array[16][6][12] <= img[7140];\
        in_img_array[16][6][13] <= img[7141];\
        in_img_array[16][6][14] <= img[7142];\
        in_img_array[16][6][15] <= img[7143];\
        in_img_array[16][6][16] <= img[7144];\
        in_img_array[16][6][17] <= img[7145];\
        in_img_array[16][7][0] <= img[7146];\
        in_img_array[16][7][1] <= img[7147];\
        in_img_array[16][7][2] <= img[7148];\
        in_img_array[16][7][3] <= img[7149];\
        in_img_array[16][7][4] <= img[7150];\
        in_img_array[16][7][5] <= img[7151];\
        in_img_array[16][7][6] <= img[7152];\
        in_img_array[16][7][7] <= img[7153];\
        in_img_array[16][7][8] <= img[7154];\
        in_img_array[16][7][9] <= img[7155];\
        in_img_array[16][7][10] <= img[7156];\
        in_img_array[16][7][11] <= img[7157];\
        in_img_array[16][7][12] <= img[7158];\
        in_img_array[16][7][13] <= img[7159];\
        in_img_array[16][7][14] <= img[7160];\
        in_img_array[16][7][15] <= img[7161];\
        in_img_array[16][7][16] <= img[7162];\
        in_img_array[16][7][17] <= img[7163];\
        in_img_array[16][8][0] <= img[7164];\
        in_img_array[16][8][1] <= img[7165];\
        in_img_array[16][8][2] <= img[7166];\
        in_img_array[16][8][3] <= img[7167];\
        in_img_array[16][8][4] <= img[7168];\
        in_img_array[16][8][5] <= img[7169];\
        in_img_array[16][8][6] <= img[7170];\
        in_img_array[16][8][7] <= img[7171];\
        in_img_array[16][8][8] <= img[7172];\
        in_img_array[16][8][9] <= img[7173];\
        in_img_array[16][8][10] <= img[7174];\
        in_img_array[16][8][11] <= img[7175];\
        in_img_array[16][8][12] <= img[7176];\
        in_img_array[16][8][13] <= img[7177];\
        in_img_array[16][8][14] <= img[7178];\
        in_img_array[16][8][15] <= img[7179];\
        in_img_array[16][8][16] <= img[7180];\
        in_img_array[16][8][17] <= img[7181];\
        in_img_array[16][9][0] <= img[7182];\
        in_img_array[16][9][1] <= img[7183];\
        in_img_array[16][9][2] <= img[7184];\
        in_img_array[16][9][3] <= img[7185];\
        in_img_array[16][9][4] <= img[7186];\
        in_img_array[16][9][5] <= img[7187];\
        in_img_array[16][9][6] <= img[7188];\
        in_img_array[16][9][7] <= img[7189];\
        in_img_array[16][9][8] <= img[7190];\
        in_img_array[16][9][9] <= img[7191];\
        in_img_array[16][9][10] <= img[7192];\
        in_img_array[16][9][11] <= img[7193];\
        in_img_array[16][9][12] <= img[7194];\
        in_img_array[16][9][13] <= img[7195];\
        in_img_array[16][9][14] <= img[7196];\
        in_img_array[16][9][15] <= img[7197];\
        in_img_array[16][9][16] <= img[7198];\
        in_img_array[16][9][17] <= img[7199];\
        in_img_array[16][10][0] <= img[7200];\
        in_img_array[16][10][1] <= img[7201];\
        in_img_array[16][10][2] <= img[7202];\
        in_img_array[16][10][3] <= img[7203];\
        in_img_array[16][10][4] <= img[7204];\
        in_img_array[16][10][5] <= img[7205];\
        in_img_array[16][10][6] <= img[7206];\
        in_img_array[16][10][7] <= img[7207];\
        in_img_array[16][10][8] <= img[7208];\
        in_img_array[16][10][9] <= img[7209];\
        in_img_array[16][10][10] <= img[7210];\
        in_img_array[16][10][11] <= img[7211];\
        in_img_array[16][10][12] <= img[7212];\
        in_img_array[16][10][13] <= img[7213];\
        in_img_array[16][10][14] <= img[7214];\
        in_img_array[16][10][15] <= img[7215];\
        in_img_array[16][10][16] <= img[7216];\
        in_img_array[16][10][17] <= img[7217];\
        in_img_array[16][11][0] <= img[7218];\
        in_img_array[16][11][1] <= img[7219];\
        in_img_array[16][11][2] <= img[7220];\
        in_img_array[16][11][3] <= img[7221];\
        in_img_array[16][11][4] <= img[7222];\
        in_img_array[16][11][5] <= img[7223];\
        in_img_array[16][11][6] <= img[7224];\
        in_img_array[16][11][7] <= img[7225];\
        in_img_array[16][11][8] <= img[7226];\
        in_img_array[16][11][9] <= img[7227];\
        in_img_array[16][11][10] <= img[7228];\
        in_img_array[16][11][11] <= img[7229];\
        in_img_array[16][11][12] <= img[7230];\
        in_img_array[16][11][13] <= img[7231];\
        in_img_array[16][11][14] <= img[7232];\
        in_img_array[16][11][15] <= img[7233];\
        in_img_array[16][11][16] <= img[7234];\
        in_img_array[16][11][17] <= img[7235];\
        in_img_array[16][12][0] <= img[7236];\
        in_img_array[16][12][1] <= img[7237];\
        in_img_array[16][12][2] <= img[7238];\
        in_img_array[16][12][3] <= img[7239];\
        in_img_array[16][12][4] <= img[7240];\
        in_img_array[16][12][5] <= img[7241];\
        in_img_array[16][12][6] <= img[7242];\
        in_img_array[16][12][7] <= img[7243];\
        in_img_array[16][12][8] <= img[7244];\
        in_img_array[16][12][9] <= img[7245];\
        in_img_array[16][12][10] <= img[7246];\
        in_img_array[16][12][11] <= img[7247];\
        in_img_array[16][12][12] <= img[7248];\
        in_img_array[16][12][13] <= img[7249];\
        in_img_array[16][12][14] <= img[7250];\
        in_img_array[16][12][15] <= img[7251];\
        in_img_array[16][12][16] <= img[7252];\
        in_img_array[16][12][17] <= img[7253];\
        in_img_array[16][13][0] <= img[7254];\
        in_img_array[16][13][1] <= img[7255];\
        in_img_array[16][13][2] <= img[7256];\
        in_img_array[16][13][3] <= img[7257];\
        in_img_array[16][13][4] <= img[7258];\
        in_img_array[16][13][5] <= img[7259];\
        in_img_array[16][13][6] <= img[7260];\
        in_img_array[16][13][7] <= img[7261];\
        in_img_array[16][13][8] <= img[7262];\
        in_img_array[16][13][9] <= img[7263];\
        in_img_array[16][13][10] <= img[7264];\
        in_img_array[16][13][11] <= img[7265];\
        in_img_array[16][13][12] <= img[7266];\
        in_img_array[16][13][13] <= img[7267];\
        in_img_array[16][13][14] <= img[7268];\
        in_img_array[16][13][15] <= img[7269];\
        in_img_array[16][13][16] <= img[7270];\
        in_img_array[16][13][17] <= img[7271];\
        in_img_array[16][14][0] <= img[7272];\
        in_img_array[16][14][1] <= img[7273];\
        in_img_array[16][14][2] <= img[7274];\
        in_img_array[16][14][3] <= img[7275];\
        in_img_array[16][14][4] <= img[7276];\
        in_img_array[16][14][5] <= img[7277];\
        in_img_array[16][14][6] <= img[7278];\
        in_img_array[16][14][7] <= img[7279];\
        in_img_array[16][14][8] <= img[7280];\
        in_img_array[16][14][9] <= img[7281];\
        in_img_array[16][14][10] <= img[7282];\
        in_img_array[16][14][11] <= img[7283];\
        in_img_array[16][14][12] <= img[7284];\
        in_img_array[16][14][13] <= img[7285];\
        in_img_array[16][14][14] <= img[7286];\
        in_img_array[16][14][15] <= img[7287];\
        in_img_array[16][14][16] <= img[7288];\
        in_img_array[16][14][17] <= img[7289];\
        in_img_array[16][15][0] <= img[7290];\
        in_img_array[16][15][1] <= img[7291];\
        in_img_array[16][15][2] <= img[7292];\
        in_img_array[16][15][3] <= img[7293];\
        in_img_array[16][15][4] <= img[7294];\
        in_img_array[16][15][5] <= img[7295];\
        in_img_array[16][15][6] <= img[7296];\
        in_img_array[16][15][7] <= img[7297];\
        in_img_array[16][15][8] <= img[7298];\
        in_img_array[16][15][9] <= img[7299];\
        in_img_array[16][15][10] <= img[7300];\
        in_img_array[16][15][11] <= img[7301];\
        in_img_array[16][15][12] <= img[7302];\
        in_img_array[16][15][13] <= img[7303];\
        in_img_array[16][15][14] <= img[7304];\
        in_img_array[16][15][15] <= img[7305];\
        in_img_array[16][15][16] <= img[7306];\
        in_img_array[16][15][17] <= img[7307];\
        in_img_array[16][16][0] <= img[7308];\
        in_img_array[16][16][1] <= img[7309];\
        in_img_array[16][16][2] <= img[7310];\
        in_img_array[16][16][3] <= img[7311];\
        in_img_array[16][16][4] <= img[7312];\
        in_img_array[16][16][5] <= img[7313];\
        in_img_array[16][16][6] <= img[7314];\
        in_img_array[16][16][7] <= img[7315];\
        in_img_array[16][16][8] <= img[7316];\
        in_img_array[16][16][9] <= img[7317];\
        in_img_array[16][16][10] <= img[7318];\
        in_img_array[16][16][11] <= img[7319];\
        in_img_array[16][16][12] <= img[7320];\
        in_img_array[16][16][13] <= img[7321];\
        in_img_array[16][16][14] <= img[7322];\
        in_img_array[16][16][15] <= img[7323];\
        in_img_array[16][16][16] <= img[7324];\
        in_img_array[16][16][17] <= img[7325];\
        in_img_array[16][17][0] <= img[7326];\
        in_img_array[16][17][1] <= img[7327];\
        in_img_array[16][17][2] <= img[7328];\
        in_img_array[16][17][3] <= img[7329];\
        in_img_array[16][17][4] <= img[7330];\
        in_img_array[16][17][5] <= img[7331];\
        in_img_array[16][17][6] <= img[7332];\
        in_img_array[16][17][7] <= img[7333];\
        in_img_array[16][17][8] <= img[7334];\
        in_img_array[16][17][9] <= img[7335];\
        in_img_array[16][17][10] <= img[7336];\
        in_img_array[16][17][11] <= img[7337];\
        in_img_array[16][17][12] <= img[7338];\
        in_img_array[16][17][13] <= img[7339];\
        in_img_array[16][17][14] <= img[7340];\
        in_img_array[16][17][15] <= img[7341];\
        in_img_array[16][17][16] <= img[7342];\
        in_img_array[16][17][17] <= img[7343];\
        in_img_array[16][18][0] <= img[7344];\
        in_img_array[16][18][1] <= img[7345];\
        in_img_array[16][18][2] <= img[7346];\
        in_img_array[16][18][3] <= img[7347];\
        in_img_array[16][18][4] <= img[7348];\
        in_img_array[16][18][5] <= img[7349];\
        in_img_array[16][18][6] <= img[7350];\
        in_img_array[16][18][7] <= img[7351];\
        in_img_array[16][18][8] <= img[7352];\
        in_img_array[16][18][9] <= img[7353];\
        in_img_array[16][18][10] <= img[7354];\
        in_img_array[16][18][11] <= img[7355];\
        in_img_array[16][18][12] <= img[7356];\
        in_img_array[16][18][13] <= img[7357];\
        in_img_array[16][18][14] <= img[7358];\
        in_img_array[16][18][15] <= img[7359];\
        in_img_array[16][18][16] <= img[7360];\
        in_img_array[16][18][17] <= img[7361];\
        in_img_array[16][19][0] <= img[7362];\
        in_img_array[16][19][1] <= img[7363];\
        in_img_array[16][19][2] <= img[7364];\
        in_img_array[16][19][3] <= img[7365];\
        in_img_array[16][19][4] <= img[7366];\
        in_img_array[16][19][5] <= img[7367];\
        in_img_array[16][19][6] <= img[7368];\
        in_img_array[16][19][7] <= img[7369];\
        in_img_array[16][19][8] <= img[7370];\
        in_img_array[16][19][9] <= img[7371];\
        in_img_array[16][19][10] <= img[7372];\
        in_img_array[16][19][11] <= img[7373];\
        in_img_array[16][19][12] <= img[7374];\
        in_img_array[16][19][13] <= img[7375];\
        in_img_array[16][19][14] <= img[7376];\
        in_img_array[16][19][15] <= img[7377];\
        in_img_array[16][19][16] <= img[7378];\
        in_img_array[16][19][17] <= img[7379];\
        in_img_array[16][20][0] <= img[7380];\
        in_img_array[16][20][1] <= img[7381];\
        in_img_array[16][20][2] <= img[7382];\
        in_img_array[16][20][3] <= img[7383];\
        in_img_array[16][20][4] <= img[7384];\
        in_img_array[16][20][5] <= img[7385];\
        in_img_array[16][20][6] <= img[7386];\
        in_img_array[16][20][7] <= img[7387];\
        in_img_array[16][20][8] <= img[7388];\
        in_img_array[16][20][9] <= img[7389];\
        in_img_array[16][20][10] <= img[7390];\
        in_img_array[16][20][11] <= img[7391];\
        in_img_array[16][20][12] <= img[7392];\
        in_img_array[16][20][13] <= img[7393];\
        in_img_array[16][20][14] <= img[7394];\
        in_img_array[16][20][15] <= img[7395];\
        in_img_array[16][20][16] <= img[7396];\
        in_img_array[16][20][17] <= img[7397];\
        in_img_array[16][21][0] <= img[7398];\
        in_img_array[16][21][1] <= img[7399];\
        in_img_array[16][21][2] <= img[7400];\
        in_img_array[16][21][3] <= img[7401];\
        in_img_array[16][21][4] <= img[7402];\
        in_img_array[16][21][5] <= img[7403];\
        in_img_array[16][21][6] <= img[7404];\
        in_img_array[16][21][7] <= img[7405];\
        in_img_array[16][21][8] <= img[7406];\
        in_img_array[16][21][9] <= img[7407];\
        in_img_array[16][21][10] <= img[7408];\
        in_img_array[16][21][11] <= img[7409];\
        in_img_array[16][21][12] <= img[7410];\
        in_img_array[16][21][13] <= img[7411];\
        in_img_array[16][21][14] <= img[7412];\
        in_img_array[16][21][15] <= img[7413];\
        in_img_array[16][21][16] <= img[7414];\
        in_img_array[16][21][17] <= img[7415];\
        in_img_array[16][22][0] <= img[7416];\
        in_img_array[16][22][1] <= img[7417];\
        in_img_array[16][22][2] <= img[7418];\
        in_img_array[16][22][3] <= img[7419];\
        in_img_array[16][22][4] <= img[7420];\
        in_img_array[16][22][5] <= img[7421];\
        in_img_array[16][22][6] <= img[7422];\
        in_img_array[16][22][7] <= img[7423];\
        in_img_array[16][22][8] <= img[7424];\
        in_img_array[16][22][9] <= img[7425];\
        in_img_array[16][22][10] <= img[7426];\
        in_img_array[16][22][11] <= img[7427];\
        in_img_array[16][22][12] <= img[7428];\
        in_img_array[16][22][13] <= img[7429];\
        in_img_array[16][22][14] <= img[7430];\
        in_img_array[16][22][15] <= img[7431];\
        in_img_array[16][22][16] <= img[7432];\
        in_img_array[16][22][17] <= img[7433];\
        in_img_array[16][23][0] <= img[7434];\
        in_img_array[16][23][1] <= img[7435];\
        in_img_array[16][23][2] <= img[7436];\
        in_img_array[16][23][3] <= img[7437];\
        in_img_array[16][23][4] <= img[7438];\
        in_img_array[16][23][5] <= img[7439];\
        in_img_array[16][23][6] <= img[7440];\
        in_img_array[16][23][7] <= img[7441];\
        in_img_array[16][23][8] <= img[7442];\
        in_img_array[16][23][9] <= img[7443];\
        in_img_array[16][23][10] <= img[7444];\
        in_img_array[16][23][11] <= img[7445];\
        in_img_array[16][23][12] <= img[7446];\
        in_img_array[16][23][13] <= img[7447];\
        in_img_array[16][23][14] <= img[7448];\
        in_img_array[16][23][15] <= img[7449];\
        in_img_array[16][23][16] <= img[7450];\
        in_img_array[16][23][17] <= img[7451];\
        in_img_array[16][24][0] <= img[7452];\
        in_img_array[16][24][1] <= img[7453];\
        in_img_array[16][24][2] <= img[7454];\
        in_img_array[16][24][3] <= img[7455];\
        in_img_array[16][24][4] <= img[7456];\
        in_img_array[16][24][5] <= img[7457];\
        in_img_array[16][24][6] <= img[7458];\
        in_img_array[16][24][7] <= img[7459];\
        in_img_array[16][24][8] <= img[7460];\
        in_img_array[16][24][9] <= img[7461];\
        in_img_array[16][24][10] <= img[7462];\
        in_img_array[16][24][11] <= img[7463];\
        in_img_array[16][24][12] <= img[7464];\
        in_img_array[16][24][13] <= img[7465];\
        in_img_array[16][24][14] <= img[7466];\
        in_img_array[16][24][15] <= img[7467];\
        in_img_array[16][24][16] <= img[7468];\
        in_img_array[16][24][17] <= img[7469];\
        in_img_array[16][25][0] <= img[7470];\
        in_img_array[16][25][1] <= img[7471];\
        in_img_array[16][25][2] <= img[7472];\
        in_img_array[16][25][3] <= img[7473];\
        in_img_array[16][25][4] <= img[7474];\
        in_img_array[16][25][5] <= img[7475];\
        in_img_array[16][25][6] <= img[7476];\
        in_img_array[16][25][7] <= img[7477];\
        in_img_array[16][25][8] <= img[7478];\
        in_img_array[16][25][9] <= img[7479];\
        in_img_array[16][25][10] <= img[7480];\
        in_img_array[16][25][11] <= img[7481];\
        in_img_array[16][25][12] <= img[7482];\
        in_img_array[16][25][13] <= img[7483];\
        in_img_array[16][25][14] <= img[7484];\
        in_img_array[16][25][15] <= img[7485];\
        in_img_array[16][25][16] <= img[7486];\
        in_img_array[16][25][17] <= img[7487];\
        in_img_array[16][26][0] <= img[7488];\
        in_img_array[16][26][1] <= img[7489];\
        in_img_array[16][26][2] <= img[7490];\
        in_img_array[16][26][3] <= img[7491];\
        in_img_array[16][26][4] <= img[7492];\
        in_img_array[16][26][5] <= img[7493];\
        in_img_array[16][26][6] <= img[7494];\
        in_img_array[16][26][7] <= img[7495];\
        in_img_array[16][26][8] <= img[7496];\
        in_img_array[16][26][9] <= img[7497];\
        in_img_array[16][26][10] <= img[7498];\
        in_img_array[16][26][11] <= img[7499];\
        in_img_array[16][26][12] <= img[7500];\
        in_img_array[16][26][13] <= img[7501];\
        in_img_array[16][26][14] <= img[7502];\
        in_img_array[16][26][15] <= img[7503];\
        in_img_array[16][26][16] <= img[7504];\
        in_img_array[16][26][17] <= img[7505];\
        in_img_array[16][27][0] <= img[7506];\
        in_img_array[16][27][1] <= img[7507];\
        in_img_array[16][27][2] <= img[7508];\
        in_img_array[16][27][3] <= img[7509];\
        in_img_array[16][27][4] <= img[7510];\
        in_img_array[16][27][5] <= img[7511];\
        in_img_array[16][27][6] <= img[7512];\
        in_img_array[16][27][7] <= img[7513];\
        in_img_array[16][27][8] <= img[7514];\
        in_img_array[16][27][9] <= img[7515];\
        in_img_array[16][27][10] <= img[7516];\
        in_img_array[16][27][11] <= img[7517];\
        in_img_array[16][27][12] <= img[7518];\
        in_img_array[16][27][13] <= img[7519];\
        in_img_array[16][27][14] <= img[7520];\
        in_img_array[16][27][15] <= img[7521];\
        in_img_array[16][27][16] <= img[7522];\
        in_img_array[16][27][17] <= img[7523];\
        in_img_array[16][28][0] <= img[7524];\
        in_img_array[16][28][1] <= img[7525];\
        in_img_array[16][28][2] <= img[7526];\
        in_img_array[16][28][3] <= img[7527];\
        in_img_array[16][28][4] <= img[7528];\
        in_img_array[16][28][5] <= img[7529];\
        in_img_array[16][28][6] <= img[7530];\
        in_img_array[16][28][7] <= img[7531];\
        in_img_array[16][28][8] <= img[7532];\
        in_img_array[16][28][9] <= img[7533];\
        in_img_array[16][28][10] <= img[7534];\
        in_img_array[16][28][11] <= img[7535];\
        in_img_array[16][28][12] <= img[7536];\
        in_img_array[16][28][13] <= img[7537];\
        in_img_array[16][28][14] <= img[7538];\
        in_img_array[16][28][15] <= img[7539];\
        in_img_array[16][28][16] <= img[7540];\
        in_img_array[16][28][17] <= img[7541];\
        in_img_array[16][29][0] <= img[7542];\
        in_img_array[16][29][1] <= img[7543];\
        in_img_array[16][29][2] <= img[7544];\
        in_img_array[16][29][3] <= img[7545];\
        in_img_array[16][29][4] <= img[7546];\
        in_img_array[16][29][5] <= img[7547];\
        in_img_array[16][29][6] <= img[7548];\
        in_img_array[16][29][7] <= img[7549];\
        in_img_array[16][29][8] <= img[7550];\
        in_img_array[16][29][9] <= img[7551];\
        in_img_array[16][29][10] <= img[7552];\
        in_img_array[16][29][11] <= img[7553];\
        in_img_array[16][29][12] <= img[7554];\
        in_img_array[16][29][13] <= img[7555];\
        in_img_array[16][29][14] <= img[7556];\
        in_img_array[16][29][15] <= img[7557];\
        in_img_array[16][29][16] <= img[7558];\
        in_img_array[16][29][17] <= img[7559];\
        in_img_array[17][2][0] <= img[7560];\
        in_img_array[17][2][1] <= img[7561];\
        in_img_array[17][2][2] <= img[7562];\
        in_img_array[17][2][3] <= img[7563];\
        in_img_array[17][2][4] <= img[7564];\
        in_img_array[17][2][5] <= img[7565];\
        in_img_array[17][2][6] <= img[7566];\
        in_img_array[17][2][7] <= img[7567];\
        in_img_array[17][2][8] <= img[7568];\
        in_img_array[17][2][9] <= img[7569];\
        in_img_array[17][2][10] <= img[7570];\
        in_img_array[17][2][11] <= img[7571];\
        in_img_array[17][2][12] <= img[7572];\
        in_img_array[17][2][13] <= img[7573];\
        in_img_array[17][2][14] <= img[7574];\
        in_img_array[17][2][15] <= img[7575];\
        in_img_array[17][2][16] <= img[7576];\
        in_img_array[17][2][17] <= img[7577];\
        in_img_array[17][3][0] <= img[7578];\
        in_img_array[17][3][1] <= img[7579];\
        in_img_array[17][3][2] <= img[7580];\
        in_img_array[17][3][3] <= img[7581];\
        in_img_array[17][3][4] <= img[7582];\
        in_img_array[17][3][5] <= img[7583];\
        in_img_array[17][3][6] <= img[7584];\
        in_img_array[17][3][7] <= img[7585];\
        in_img_array[17][3][8] <= img[7586];\
        in_img_array[17][3][9] <= img[7587];\
        in_img_array[17][3][10] <= img[7588];\
        in_img_array[17][3][11] <= img[7589];\
        in_img_array[17][3][12] <= img[7590];\
        in_img_array[17][3][13] <= img[7591];\
        in_img_array[17][3][14] <= img[7592];\
        in_img_array[17][3][15] <= img[7593];\
        in_img_array[17][3][16] <= img[7594];\
        in_img_array[17][3][17] <= img[7595];\
        in_img_array[17][4][0] <= img[7596];\
        in_img_array[17][4][1] <= img[7597];\
        in_img_array[17][4][2] <= img[7598];\
        in_img_array[17][4][3] <= img[7599];\
        in_img_array[17][4][4] <= img[7600];\
        in_img_array[17][4][5] <= img[7601];\
        in_img_array[17][4][6] <= img[7602];\
        in_img_array[17][4][7] <= img[7603];\
        in_img_array[17][4][8] <= img[7604];\
        in_img_array[17][4][9] <= img[7605];\
        in_img_array[17][4][10] <= img[7606];\
        in_img_array[17][4][11] <= img[7607];\
        in_img_array[17][4][12] <= img[7608];\
        in_img_array[17][4][13] <= img[7609];\
        in_img_array[17][4][14] <= img[7610];\
        in_img_array[17][4][15] <= img[7611];\
        in_img_array[17][4][16] <= img[7612];\
        in_img_array[17][4][17] <= img[7613];\
        in_img_array[17][5][0] <= img[7614];\
        in_img_array[17][5][1] <= img[7615];\
        in_img_array[17][5][2] <= img[7616];\
        in_img_array[17][5][3] <= img[7617];\
        in_img_array[17][5][4] <= img[7618];\
        in_img_array[17][5][5] <= img[7619];\
        in_img_array[17][5][6] <= img[7620];\
        in_img_array[17][5][7] <= img[7621];\
        in_img_array[17][5][8] <= img[7622];\
        in_img_array[17][5][9] <= img[7623];\
        in_img_array[17][5][10] <= img[7624];\
        in_img_array[17][5][11] <= img[7625];\
        in_img_array[17][5][12] <= img[7626];\
        in_img_array[17][5][13] <= img[7627];\
        in_img_array[17][5][14] <= img[7628];\
        in_img_array[17][5][15] <= img[7629];\
        in_img_array[17][5][16] <= img[7630];\
        in_img_array[17][5][17] <= img[7631];\
        in_img_array[17][6][0] <= img[7632];\
        in_img_array[17][6][1] <= img[7633];\
        in_img_array[17][6][2] <= img[7634];\
        in_img_array[17][6][3] <= img[7635];\
        in_img_array[17][6][4] <= img[7636];\
        in_img_array[17][6][5] <= img[7637];\
        in_img_array[17][6][6] <= img[7638];\
        in_img_array[17][6][7] <= img[7639];\
        in_img_array[17][6][8] <= img[7640];\
        in_img_array[17][6][9] <= img[7641];\
        in_img_array[17][6][10] <= img[7642];\
        in_img_array[17][6][11] <= img[7643];\
        in_img_array[17][6][12] <= img[7644];\
        in_img_array[17][6][13] <= img[7645];\
        in_img_array[17][6][14] <= img[7646];\
        in_img_array[17][6][15] <= img[7647];\
        in_img_array[17][6][16] <= img[7648];\
        in_img_array[17][6][17] <= img[7649];\
        in_img_array[17][7][0] <= img[7650];\
        in_img_array[17][7][1] <= img[7651];\
        in_img_array[17][7][2] <= img[7652];\
        in_img_array[17][7][3] <= img[7653];\
        in_img_array[17][7][4] <= img[7654];\
        in_img_array[17][7][5] <= img[7655];\
        in_img_array[17][7][6] <= img[7656];\
        in_img_array[17][7][7] <= img[7657];\
        in_img_array[17][7][8] <= img[7658];\
        in_img_array[17][7][9] <= img[7659];\
        in_img_array[17][7][10] <= img[7660];\
        in_img_array[17][7][11] <= img[7661];\
        in_img_array[17][7][12] <= img[7662];\
        in_img_array[17][7][13] <= img[7663];\
        in_img_array[17][7][14] <= img[7664];\
        in_img_array[17][7][15] <= img[7665];\
        in_img_array[17][7][16] <= img[7666];\
        in_img_array[17][7][17] <= img[7667];\
        in_img_array[17][8][0] <= img[7668];\
        in_img_array[17][8][1] <= img[7669];\
        in_img_array[17][8][2] <= img[7670];\
        in_img_array[17][8][3] <= img[7671];\
        in_img_array[17][8][4] <= img[7672];\
        in_img_array[17][8][5] <= img[7673];\
        in_img_array[17][8][6] <= img[7674];\
        in_img_array[17][8][7] <= img[7675];\
        in_img_array[17][8][8] <= img[7676];\
        in_img_array[17][8][9] <= img[7677];\
        in_img_array[17][8][10] <= img[7678];\
        in_img_array[17][8][11] <= img[7679];\
        in_img_array[17][8][12] <= img[7680];\
        in_img_array[17][8][13] <= img[7681];\
        in_img_array[17][8][14] <= img[7682];\
        in_img_array[17][8][15] <= img[7683];\
        in_img_array[17][8][16] <= img[7684];\
        in_img_array[17][8][17] <= img[7685];\
        in_img_array[17][9][0] <= img[7686];\
        in_img_array[17][9][1] <= img[7687];\
        in_img_array[17][9][2] <= img[7688];\
        in_img_array[17][9][3] <= img[7689];\
        in_img_array[17][9][4] <= img[7690];\
        in_img_array[17][9][5] <= img[7691];\
        in_img_array[17][9][6] <= img[7692];\
        in_img_array[17][9][7] <= img[7693];\
        in_img_array[17][9][8] <= img[7694];\
        in_img_array[17][9][9] <= img[7695];\
        in_img_array[17][9][10] <= img[7696];\
        in_img_array[17][9][11] <= img[7697];\
        in_img_array[17][9][12] <= img[7698];\
        in_img_array[17][9][13] <= img[7699];\
        in_img_array[17][9][14] <= img[7700];\
        in_img_array[17][9][15] <= img[7701];\
        in_img_array[17][9][16] <= img[7702];\
        in_img_array[17][9][17] <= img[7703];\
        in_img_array[17][10][0] <= img[7704];\
        in_img_array[17][10][1] <= img[7705];\
        in_img_array[17][10][2] <= img[7706];\
        in_img_array[17][10][3] <= img[7707];\
        in_img_array[17][10][4] <= img[7708];\
        in_img_array[17][10][5] <= img[7709];\
        in_img_array[17][10][6] <= img[7710];\
        in_img_array[17][10][7] <= img[7711];\
        in_img_array[17][10][8] <= img[7712];\
        in_img_array[17][10][9] <= img[7713];\
        in_img_array[17][10][10] <= img[7714];\
        in_img_array[17][10][11] <= img[7715];\
        in_img_array[17][10][12] <= img[7716];\
        in_img_array[17][10][13] <= img[7717];\
        in_img_array[17][10][14] <= img[7718];\
        in_img_array[17][10][15] <= img[7719];\
        in_img_array[17][10][16] <= img[7720];\
        in_img_array[17][10][17] <= img[7721];\
        in_img_array[17][11][0] <= img[7722];\
        in_img_array[17][11][1] <= img[7723];\
        in_img_array[17][11][2] <= img[7724];\
        in_img_array[17][11][3] <= img[7725];\
        in_img_array[17][11][4] <= img[7726];\
        in_img_array[17][11][5] <= img[7727];\
        in_img_array[17][11][6] <= img[7728];\
        in_img_array[17][11][7] <= img[7729];\
        in_img_array[17][11][8] <= img[7730];\
        in_img_array[17][11][9] <= img[7731];\
        in_img_array[17][11][10] <= img[7732];\
        in_img_array[17][11][11] <= img[7733];\
        in_img_array[17][11][12] <= img[7734];\
        in_img_array[17][11][13] <= img[7735];\
        in_img_array[17][11][14] <= img[7736];\
        in_img_array[17][11][15] <= img[7737];\
        in_img_array[17][11][16] <= img[7738];\
        in_img_array[17][11][17] <= img[7739];\
        in_img_array[17][12][0] <= img[7740];\
        in_img_array[17][12][1] <= img[7741];\
        in_img_array[17][12][2] <= img[7742];\
        in_img_array[17][12][3] <= img[7743];\
        in_img_array[17][12][4] <= img[7744];\
        in_img_array[17][12][5] <= img[7745];\
        in_img_array[17][12][6] <= img[7746];\
        in_img_array[17][12][7] <= img[7747];\
        in_img_array[17][12][8] <= img[7748];\
        in_img_array[17][12][9] <= img[7749];\
        in_img_array[17][12][10] <= img[7750];\
        in_img_array[17][12][11] <= img[7751];\
        in_img_array[17][12][12] <= img[7752];\
        in_img_array[17][12][13] <= img[7753];\
        in_img_array[17][12][14] <= img[7754];\
        in_img_array[17][12][15] <= img[7755];\
        in_img_array[17][12][16] <= img[7756];\
        in_img_array[17][12][17] <= img[7757];\
        in_img_array[17][13][0] <= img[7758];\
        in_img_array[17][13][1] <= img[7759];\
        in_img_array[17][13][2] <= img[7760];\
        in_img_array[17][13][3] <= img[7761];\
        in_img_array[17][13][4] <= img[7762];\
        in_img_array[17][13][5] <= img[7763];\
        in_img_array[17][13][6] <= img[7764];\
        in_img_array[17][13][7] <= img[7765];\
        in_img_array[17][13][8] <= img[7766];\
        in_img_array[17][13][9] <= img[7767];\
        in_img_array[17][13][10] <= img[7768];\
        in_img_array[17][13][11] <= img[7769];\
        in_img_array[17][13][12] <= img[7770];\
        in_img_array[17][13][13] <= img[7771];\
        in_img_array[17][13][14] <= img[7772];\
        in_img_array[17][13][15] <= img[7773];\
        in_img_array[17][13][16] <= img[7774];\
        in_img_array[17][13][17] <= img[7775];\
        in_img_array[17][14][0] <= img[7776];\
        in_img_array[17][14][1] <= img[7777];\
        in_img_array[17][14][2] <= img[7778];\
        in_img_array[17][14][3] <= img[7779];\
        in_img_array[17][14][4] <= img[7780];\
        in_img_array[17][14][5] <= img[7781];\
        in_img_array[17][14][6] <= img[7782];\
        in_img_array[17][14][7] <= img[7783];\
        in_img_array[17][14][8] <= img[7784];\
        in_img_array[17][14][9] <= img[7785];\
        in_img_array[17][14][10] <= img[7786];\
        in_img_array[17][14][11] <= img[7787];\
        in_img_array[17][14][12] <= img[7788];\
        in_img_array[17][14][13] <= img[7789];\
        in_img_array[17][14][14] <= img[7790];\
        in_img_array[17][14][15] <= img[7791];\
        in_img_array[17][14][16] <= img[7792];\
        in_img_array[17][14][17] <= img[7793];\
        in_img_array[17][15][0] <= img[7794];\
        in_img_array[17][15][1] <= img[7795];\
        in_img_array[17][15][2] <= img[7796];\
        in_img_array[17][15][3] <= img[7797];\
        in_img_array[17][15][4] <= img[7798];\
        in_img_array[17][15][5] <= img[7799];\
        in_img_array[17][15][6] <= img[7800];\
        in_img_array[17][15][7] <= img[7801];\
        in_img_array[17][15][8] <= img[7802];\
        in_img_array[17][15][9] <= img[7803];\
        in_img_array[17][15][10] <= img[7804];\
        in_img_array[17][15][11] <= img[7805];\
        in_img_array[17][15][12] <= img[7806];\
        in_img_array[17][15][13] <= img[7807];\
        in_img_array[17][15][14] <= img[7808];\
        in_img_array[17][15][15] <= img[7809];\
        in_img_array[17][15][16] <= img[7810];\
        in_img_array[17][15][17] <= img[7811];\
        in_img_array[17][16][0] <= img[7812];\
        in_img_array[17][16][1] <= img[7813];\
        in_img_array[17][16][2] <= img[7814];\
        in_img_array[17][16][3] <= img[7815];\
        in_img_array[17][16][4] <= img[7816];\
        in_img_array[17][16][5] <= img[7817];\
        in_img_array[17][16][6] <= img[7818];\
        in_img_array[17][16][7] <= img[7819];\
        in_img_array[17][16][8] <= img[7820];\
        in_img_array[17][16][9] <= img[7821];\
        in_img_array[17][16][10] <= img[7822];\
        in_img_array[17][16][11] <= img[7823];\
        in_img_array[17][16][12] <= img[7824];\
        in_img_array[17][16][13] <= img[7825];\
        in_img_array[17][16][14] <= img[7826];\
        in_img_array[17][16][15] <= img[7827];\
        in_img_array[17][16][16] <= img[7828];\
        in_img_array[17][16][17] <= img[7829];\
        in_img_array[17][17][0] <= img[7830];\
        in_img_array[17][17][1] <= img[7831];\
        in_img_array[17][17][2] <= img[7832];\
        in_img_array[17][17][3] <= img[7833];\
        in_img_array[17][17][4] <= img[7834];\
        in_img_array[17][17][5] <= img[7835];\
        in_img_array[17][17][6] <= img[7836];\
        in_img_array[17][17][7] <= img[7837];\
        in_img_array[17][17][8] <= img[7838];\
        in_img_array[17][17][9] <= img[7839];\
        in_img_array[17][17][10] <= img[7840];\
        in_img_array[17][17][11] <= img[7841];\
        in_img_array[17][17][12] <= img[7842];\
        in_img_array[17][17][13] <= img[7843];\
        in_img_array[17][17][14] <= img[7844];\
        in_img_array[17][17][15] <= img[7845];\
        in_img_array[17][17][16] <= img[7846];\
        in_img_array[17][17][17] <= img[7847];\
        in_img_array[17][18][0] <= img[7848];\
        in_img_array[17][18][1] <= img[7849];\
        in_img_array[17][18][2] <= img[7850];\
        in_img_array[17][18][3] <= img[7851];\
        in_img_array[17][18][4] <= img[7852];\
        in_img_array[17][18][5] <= img[7853];\
        in_img_array[17][18][6] <= img[7854];\
        in_img_array[17][18][7] <= img[7855];\
        in_img_array[17][18][8] <= img[7856];\
        in_img_array[17][18][9] <= img[7857];\
        in_img_array[17][18][10] <= img[7858];\
        in_img_array[17][18][11] <= img[7859];\
        in_img_array[17][18][12] <= img[7860];\
        in_img_array[17][18][13] <= img[7861];\
        in_img_array[17][18][14] <= img[7862];\
        in_img_array[17][18][15] <= img[7863];\
        in_img_array[17][18][16] <= img[7864];\
        in_img_array[17][18][17] <= img[7865];\
        in_img_array[17][19][0] <= img[7866];\
        in_img_array[17][19][1] <= img[7867];\
        in_img_array[17][19][2] <= img[7868];\
        in_img_array[17][19][3] <= img[7869];\
        in_img_array[17][19][4] <= img[7870];\
        in_img_array[17][19][5] <= img[7871];\
        in_img_array[17][19][6] <= img[7872];\
        in_img_array[17][19][7] <= img[7873];\
        in_img_array[17][19][8] <= img[7874];\
        in_img_array[17][19][9] <= img[7875];\
        in_img_array[17][19][10] <= img[7876];\
        in_img_array[17][19][11] <= img[7877];\
        in_img_array[17][19][12] <= img[7878];\
        in_img_array[17][19][13] <= img[7879];\
        in_img_array[17][19][14] <= img[7880];\
        in_img_array[17][19][15] <= img[7881];\
        in_img_array[17][19][16] <= img[7882];\
        in_img_array[17][19][17] <= img[7883];\
        in_img_array[17][20][0] <= img[7884];\
        in_img_array[17][20][1] <= img[7885];\
        in_img_array[17][20][2] <= img[7886];\
        in_img_array[17][20][3] <= img[7887];\
        in_img_array[17][20][4] <= img[7888];\
        in_img_array[17][20][5] <= img[7889];\
        in_img_array[17][20][6] <= img[7890];\
        in_img_array[17][20][7] <= img[7891];\
        in_img_array[17][20][8] <= img[7892];\
        in_img_array[17][20][9] <= img[7893];\
        in_img_array[17][20][10] <= img[7894];\
        in_img_array[17][20][11] <= img[7895];\
        in_img_array[17][20][12] <= img[7896];\
        in_img_array[17][20][13] <= img[7897];\
        in_img_array[17][20][14] <= img[7898];\
        in_img_array[17][20][15] <= img[7899];\
        in_img_array[17][20][16] <= img[7900];\
        in_img_array[17][20][17] <= img[7901];\
        in_img_array[17][21][0] <= img[7902];\
        in_img_array[17][21][1] <= img[7903];\
        in_img_array[17][21][2] <= img[7904];\
        in_img_array[17][21][3] <= img[7905];\
        in_img_array[17][21][4] <= img[7906];\
        in_img_array[17][21][5] <= img[7907];\
        in_img_array[17][21][6] <= img[7908];\
        in_img_array[17][21][7] <= img[7909];\
        in_img_array[17][21][8] <= img[7910];\
        in_img_array[17][21][9] <= img[7911];\
        in_img_array[17][21][10] <= img[7912];\
        in_img_array[17][21][11] <= img[7913];\
        in_img_array[17][21][12] <= img[7914];\
        in_img_array[17][21][13] <= img[7915];\
        in_img_array[17][21][14] <= img[7916];\
        in_img_array[17][21][15] <= img[7917];\
        in_img_array[17][21][16] <= img[7918];\
        in_img_array[17][21][17] <= img[7919];\
        in_img_array[17][22][0] <= img[7920];\
        in_img_array[17][22][1] <= img[7921];\
        in_img_array[17][22][2] <= img[7922];\
        in_img_array[17][22][3] <= img[7923];\
        in_img_array[17][22][4] <= img[7924];\
        in_img_array[17][22][5] <= img[7925];\
        in_img_array[17][22][6] <= img[7926];\
        in_img_array[17][22][7] <= img[7927];\
        in_img_array[17][22][8] <= img[7928];\
        in_img_array[17][22][9] <= img[7929];\
        in_img_array[17][22][10] <= img[7930];\
        in_img_array[17][22][11] <= img[7931];\
        in_img_array[17][22][12] <= img[7932];\
        in_img_array[17][22][13] <= img[7933];\
        in_img_array[17][22][14] <= img[7934];\
        in_img_array[17][22][15] <= img[7935];\
        in_img_array[17][22][16] <= img[7936];\
        in_img_array[17][22][17] <= img[7937];\
        in_img_array[17][23][0] <= img[7938];\
        in_img_array[17][23][1] <= img[7939];\
        in_img_array[17][23][2] <= img[7940];\
        in_img_array[17][23][3] <= img[7941];\
        in_img_array[17][23][4] <= img[7942];\
        in_img_array[17][23][5] <= img[7943];\
        in_img_array[17][23][6] <= img[7944];\
        in_img_array[17][23][7] <= img[7945];\
        in_img_array[17][23][8] <= img[7946];\
        in_img_array[17][23][9] <= img[7947];\
        in_img_array[17][23][10] <= img[7948];\
        in_img_array[17][23][11] <= img[7949];\
        in_img_array[17][23][12] <= img[7950];\
        in_img_array[17][23][13] <= img[7951];\
        in_img_array[17][23][14] <= img[7952];\
        in_img_array[17][23][15] <= img[7953];\
        in_img_array[17][23][16] <= img[7954];\
        in_img_array[17][23][17] <= img[7955];\
        in_img_array[17][24][0] <= img[7956];\
        in_img_array[17][24][1] <= img[7957];\
        in_img_array[17][24][2] <= img[7958];\
        in_img_array[17][24][3] <= img[7959];\
        in_img_array[17][24][4] <= img[7960];\
        in_img_array[17][24][5] <= img[7961];\
        in_img_array[17][24][6] <= img[7962];\
        in_img_array[17][24][7] <= img[7963];\
        in_img_array[17][24][8] <= img[7964];\
        in_img_array[17][24][9] <= img[7965];\
        in_img_array[17][24][10] <= img[7966];\
        in_img_array[17][24][11] <= img[7967];\
        in_img_array[17][24][12] <= img[7968];\
        in_img_array[17][24][13] <= img[7969];\
        in_img_array[17][24][14] <= img[7970];\
        in_img_array[17][24][15] <= img[7971];\
        in_img_array[17][24][16] <= img[7972];\
        in_img_array[17][24][17] <= img[7973];\
        in_img_array[17][25][0] <= img[7974];\
        in_img_array[17][25][1] <= img[7975];\
        in_img_array[17][25][2] <= img[7976];\
        in_img_array[17][25][3] <= img[7977];\
        in_img_array[17][25][4] <= img[7978];\
        in_img_array[17][25][5] <= img[7979];\
        in_img_array[17][25][6] <= img[7980];\
        in_img_array[17][25][7] <= img[7981];\
        in_img_array[17][25][8] <= img[7982];\
        in_img_array[17][25][9] <= img[7983];\
        in_img_array[17][25][10] <= img[7984];\
        in_img_array[17][25][11] <= img[7985];\
        in_img_array[17][25][12] <= img[7986];\
        in_img_array[17][25][13] <= img[7987];\
        in_img_array[17][25][14] <= img[7988];\
        in_img_array[17][25][15] <= img[7989];\
        in_img_array[17][25][16] <= img[7990];\
        in_img_array[17][25][17] <= img[7991];\
        in_img_array[17][26][0] <= img[7992];\
        in_img_array[17][26][1] <= img[7993];\
        in_img_array[17][26][2] <= img[7994];\
        in_img_array[17][26][3] <= img[7995];\
        in_img_array[17][26][4] <= img[7996];\
        in_img_array[17][26][5] <= img[7997];\
        in_img_array[17][26][6] <= img[7998];\
        in_img_array[17][26][7] <= img[7999];\
        in_img_array[17][26][8] <= img[8000];\
        in_img_array[17][26][9] <= img[8001];\
        in_img_array[17][26][10] <= img[8002];\
        in_img_array[17][26][11] <= img[8003];\
        in_img_array[17][26][12] <= img[8004];\
        in_img_array[17][26][13] <= img[8005];\
        in_img_array[17][26][14] <= img[8006];\
        in_img_array[17][26][15] <= img[8007];\
        in_img_array[17][26][16] <= img[8008];\
        in_img_array[17][26][17] <= img[8009];\
        in_img_array[17][27][0] <= img[8010];\
        in_img_array[17][27][1] <= img[8011];\
        in_img_array[17][27][2] <= img[8012];\
        in_img_array[17][27][3] <= img[8013];\
        in_img_array[17][27][4] <= img[8014];\
        in_img_array[17][27][5] <= img[8015];\
        in_img_array[17][27][6] <= img[8016];\
        in_img_array[17][27][7] <= img[8017];\
        in_img_array[17][27][8] <= img[8018];\
        in_img_array[17][27][9] <= img[8019];\
        in_img_array[17][27][10] <= img[8020];\
        in_img_array[17][27][11] <= img[8021];\
        in_img_array[17][27][12] <= img[8022];\
        in_img_array[17][27][13] <= img[8023];\
        in_img_array[17][27][14] <= img[8024];\
        in_img_array[17][27][15] <= img[8025];\
        in_img_array[17][27][16] <= img[8026];\
        in_img_array[17][27][17] <= img[8027];\
        in_img_array[17][28][0] <= img[8028];\
        in_img_array[17][28][1] <= img[8029];\
        in_img_array[17][28][2] <= img[8030];\
        in_img_array[17][28][3] <= img[8031];\
        in_img_array[17][28][4] <= img[8032];\
        in_img_array[17][28][5] <= img[8033];\
        in_img_array[17][28][6] <= img[8034];\
        in_img_array[17][28][7] <= img[8035];\
        in_img_array[17][28][8] <= img[8036];\
        in_img_array[17][28][9] <= img[8037];\
        in_img_array[17][28][10] <= img[8038];\
        in_img_array[17][28][11] <= img[8039];\
        in_img_array[17][28][12] <= img[8040];\
        in_img_array[17][28][13] <= img[8041];\
        in_img_array[17][28][14] <= img[8042];\
        in_img_array[17][28][15] <= img[8043];\
        in_img_array[17][28][16] <= img[8044];\
        in_img_array[17][28][17] <= img[8045];\
        in_img_array[17][29][0] <= img[8046];\
        in_img_array[17][29][1] <= img[8047];\
        in_img_array[17][29][2] <= img[8048];\
        in_img_array[17][29][3] <= img[8049];\
        in_img_array[17][29][4] <= img[8050];\
        in_img_array[17][29][5] <= img[8051];\
        in_img_array[17][29][6] <= img[8052];\
        in_img_array[17][29][7] <= img[8053];\
        in_img_array[17][29][8] <= img[8054];\
        in_img_array[17][29][9] <= img[8055];\
        in_img_array[17][29][10] <= img[8056];\
        in_img_array[17][29][11] <= img[8057];\
        in_img_array[17][29][12] <= img[8058];\
        in_img_array[17][29][13] <= img[8059];\
        in_img_array[17][29][14] <= img[8060];\
        in_img_array[17][29][15] <= img[8061];\
        in_img_array[17][29][16] <= img[8062];\
        in_img_array[17][29][17] <= img[8063];\
        in_img_array[18][2][0] <= img[8064];\
        in_img_array[18][2][1] <= img[8065];\
        in_img_array[18][2][2] <= img[8066];\
        in_img_array[18][2][3] <= img[8067];\
        in_img_array[18][2][4] <= img[8068];\
        in_img_array[18][2][5] <= img[8069];\
        in_img_array[18][2][6] <= img[8070];\
        in_img_array[18][2][7] <= img[8071];\
        in_img_array[18][2][8] <= img[8072];\
        in_img_array[18][2][9] <= img[8073];\
        in_img_array[18][2][10] <= img[8074];\
        in_img_array[18][2][11] <= img[8075];\
        in_img_array[18][2][12] <= img[8076];\
        in_img_array[18][2][13] <= img[8077];\
        in_img_array[18][2][14] <= img[8078];\
        in_img_array[18][2][15] <= img[8079];\
        in_img_array[18][2][16] <= img[8080];\
        in_img_array[18][2][17] <= img[8081];\
        in_img_array[18][3][0] <= img[8082];\
        in_img_array[18][3][1] <= img[8083];\
        in_img_array[18][3][2] <= img[8084];\
        in_img_array[18][3][3] <= img[8085];\
        in_img_array[18][3][4] <= img[8086];\
        in_img_array[18][3][5] <= img[8087];\
        in_img_array[18][3][6] <= img[8088];\
        in_img_array[18][3][7] <= img[8089];\
        in_img_array[18][3][8] <= img[8090];\
        in_img_array[18][3][9] <= img[8091];\
        in_img_array[18][3][10] <= img[8092];\
        in_img_array[18][3][11] <= img[8093];\
        in_img_array[18][3][12] <= img[8094];\
        in_img_array[18][3][13] <= img[8095];\
        in_img_array[18][3][14] <= img[8096];\
        in_img_array[18][3][15] <= img[8097];\
        in_img_array[18][3][16] <= img[8098];\
        in_img_array[18][3][17] <= img[8099];\
        in_img_array[18][4][0] <= img[8100];\
        in_img_array[18][4][1] <= img[8101];\
        in_img_array[18][4][2] <= img[8102];\
        in_img_array[18][4][3] <= img[8103];\
        in_img_array[18][4][4] <= img[8104];\
        in_img_array[18][4][5] <= img[8105];\
        in_img_array[18][4][6] <= img[8106];\
        in_img_array[18][4][7] <= img[8107];\
        in_img_array[18][4][8] <= img[8108];\
        in_img_array[18][4][9] <= img[8109];\
        in_img_array[18][4][10] <= img[8110];\
        in_img_array[18][4][11] <= img[8111];\
        in_img_array[18][4][12] <= img[8112];\
        in_img_array[18][4][13] <= img[8113];\
        in_img_array[18][4][14] <= img[8114];\
        in_img_array[18][4][15] <= img[8115];\
        in_img_array[18][4][16] <= img[8116];\
        in_img_array[18][4][17] <= img[8117];\
        in_img_array[18][5][0] <= img[8118];\
        in_img_array[18][5][1] <= img[8119];\
        in_img_array[18][5][2] <= img[8120];\
        in_img_array[18][5][3] <= img[8121];\
        in_img_array[18][5][4] <= img[8122];\
        in_img_array[18][5][5] <= img[8123];\
        in_img_array[18][5][6] <= img[8124];\
        in_img_array[18][5][7] <= img[8125];\
        in_img_array[18][5][8] <= img[8126];\
        in_img_array[18][5][9] <= img[8127];\
        in_img_array[18][5][10] <= img[8128];\
        in_img_array[18][5][11] <= img[8129];\
        in_img_array[18][5][12] <= img[8130];\
        in_img_array[18][5][13] <= img[8131];\
        in_img_array[18][5][14] <= img[8132];\
        in_img_array[18][5][15] <= img[8133];\
        in_img_array[18][5][16] <= img[8134];\
        in_img_array[18][5][17] <= img[8135];\
        in_img_array[18][6][0] <= img[8136];\
        in_img_array[18][6][1] <= img[8137];\
        in_img_array[18][6][2] <= img[8138];\
        in_img_array[18][6][3] <= img[8139];\
        in_img_array[18][6][4] <= img[8140];\
        in_img_array[18][6][5] <= img[8141];\
        in_img_array[18][6][6] <= img[8142];\
        in_img_array[18][6][7] <= img[8143];\
        in_img_array[18][6][8] <= img[8144];\
        in_img_array[18][6][9] <= img[8145];\
        in_img_array[18][6][10] <= img[8146];\
        in_img_array[18][6][11] <= img[8147];\
        in_img_array[18][6][12] <= img[8148];\
        in_img_array[18][6][13] <= img[8149];\
        in_img_array[18][6][14] <= img[8150];\
        in_img_array[18][6][15] <= img[8151];\
        in_img_array[18][6][16] <= img[8152];\
        in_img_array[18][6][17] <= img[8153];\
        in_img_array[18][7][0] <= img[8154];\
        in_img_array[18][7][1] <= img[8155];\
        in_img_array[18][7][2] <= img[8156];\
        in_img_array[18][7][3] <= img[8157];\
        in_img_array[18][7][4] <= img[8158];\
        in_img_array[18][7][5] <= img[8159];\
        in_img_array[18][7][6] <= img[8160];\
        in_img_array[18][7][7] <= img[8161];\
        in_img_array[18][7][8] <= img[8162];\
        in_img_array[18][7][9] <= img[8163];\
        in_img_array[18][7][10] <= img[8164];\
        in_img_array[18][7][11] <= img[8165];\
        in_img_array[18][7][12] <= img[8166];\
        in_img_array[18][7][13] <= img[8167];\
        in_img_array[18][7][14] <= img[8168];\
        in_img_array[18][7][15] <= img[8169];\
        in_img_array[18][7][16] <= img[8170];\
        in_img_array[18][7][17] <= img[8171];\
        in_img_array[18][8][0] <= img[8172];\
        in_img_array[18][8][1] <= img[8173];\
        in_img_array[18][8][2] <= img[8174];\
        in_img_array[18][8][3] <= img[8175];\
        in_img_array[18][8][4] <= img[8176];\
        in_img_array[18][8][5] <= img[8177];\
        in_img_array[18][8][6] <= img[8178];\
        in_img_array[18][8][7] <= img[8179];\
        in_img_array[18][8][8] <= img[8180];\
        in_img_array[18][8][9] <= img[8181];\
        in_img_array[18][8][10] <= img[8182];\
        in_img_array[18][8][11] <= img[8183];\
        in_img_array[18][8][12] <= img[8184];\
        in_img_array[18][8][13] <= img[8185];\
        in_img_array[18][8][14] <= img[8186];\
        in_img_array[18][8][15] <= img[8187];\
        in_img_array[18][8][16] <= img[8188];\
        in_img_array[18][8][17] <= img[8189];\
        in_img_array[18][9][0] <= img[8190];\
        in_img_array[18][9][1] <= img[8191];\
        in_img_array[18][9][2] <= img[8192];\
        in_img_array[18][9][3] <= img[8193];\
        in_img_array[18][9][4] <= img[8194];\
        in_img_array[18][9][5] <= img[8195];\
        in_img_array[18][9][6] <= img[8196];\
        in_img_array[18][9][7] <= img[8197];\
        in_img_array[18][9][8] <= img[8198];\
        in_img_array[18][9][9] <= img[8199];\
        in_img_array[18][9][10] <= img[8200];\
        in_img_array[18][9][11] <= img[8201];\
        in_img_array[18][9][12] <= img[8202];\
        in_img_array[18][9][13] <= img[8203];\
        in_img_array[18][9][14] <= img[8204];\
        in_img_array[18][9][15] <= img[8205];\
        in_img_array[18][9][16] <= img[8206];\
        in_img_array[18][9][17] <= img[8207];\
        in_img_array[18][10][0] <= img[8208];\
        in_img_array[18][10][1] <= img[8209];\
        in_img_array[18][10][2] <= img[8210];\
        in_img_array[18][10][3] <= img[8211];\
        in_img_array[18][10][4] <= img[8212];\
        in_img_array[18][10][5] <= img[8213];\
        in_img_array[18][10][6] <= img[8214];\
        in_img_array[18][10][7] <= img[8215];\
        in_img_array[18][10][8] <= img[8216];\
        in_img_array[18][10][9] <= img[8217];\
        in_img_array[18][10][10] <= img[8218];\
        in_img_array[18][10][11] <= img[8219];\
        in_img_array[18][10][12] <= img[8220];\
        in_img_array[18][10][13] <= img[8221];\
        in_img_array[18][10][14] <= img[8222];\
        in_img_array[18][10][15] <= img[8223];\
        in_img_array[18][10][16] <= img[8224];\
        in_img_array[18][10][17] <= img[8225];\
        in_img_array[18][11][0] <= img[8226];\
        in_img_array[18][11][1] <= img[8227];\
        in_img_array[18][11][2] <= img[8228];\
        in_img_array[18][11][3] <= img[8229];\
        in_img_array[18][11][4] <= img[8230];\
        in_img_array[18][11][5] <= img[8231];\
        in_img_array[18][11][6] <= img[8232];\
        in_img_array[18][11][7] <= img[8233];\
        in_img_array[18][11][8] <= img[8234];\
        in_img_array[18][11][9] <= img[8235];\
        in_img_array[18][11][10] <= img[8236];\
        in_img_array[18][11][11] <= img[8237];\
        in_img_array[18][11][12] <= img[8238];\
        in_img_array[18][11][13] <= img[8239];\
        in_img_array[18][11][14] <= img[8240];\
        in_img_array[18][11][15] <= img[8241];\
        in_img_array[18][11][16] <= img[8242];\
        in_img_array[18][11][17] <= img[8243];\
        in_img_array[18][12][0] <= img[8244];\
        in_img_array[18][12][1] <= img[8245];\
        in_img_array[18][12][2] <= img[8246];\
        in_img_array[18][12][3] <= img[8247];\
        in_img_array[18][12][4] <= img[8248];\
        in_img_array[18][12][5] <= img[8249];\
        in_img_array[18][12][6] <= img[8250];\
        in_img_array[18][12][7] <= img[8251];\
        in_img_array[18][12][8] <= img[8252];\
        in_img_array[18][12][9] <= img[8253];\
        in_img_array[18][12][10] <= img[8254];\
        in_img_array[18][12][11] <= img[8255];\
        in_img_array[18][12][12] <= img[8256];\
        in_img_array[18][12][13] <= img[8257];\
        in_img_array[18][12][14] <= img[8258];\
        in_img_array[18][12][15] <= img[8259];\
        in_img_array[18][12][16] <= img[8260];\
        in_img_array[18][12][17] <= img[8261];\
        in_img_array[18][13][0] <= img[8262];\
        in_img_array[18][13][1] <= img[8263];\
        in_img_array[18][13][2] <= img[8264];\
        in_img_array[18][13][3] <= img[8265];\
        in_img_array[18][13][4] <= img[8266];\
        in_img_array[18][13][5] <= img[8267];\
        in_img_array[18][13][6] <= img[8268];\
        in_img_array[18][13][7] <= img[8269];\
        in_img_array[18][13][8] <= img[8270];\
        in_img_array[18][13][9] <= img[8271];\
        in_img_array[18][13][10] <= img[8272];\
        in_img_array[18][13][11] <= img[8273];\
        in_img_array[18][13][12] <= img[8274];\
        in_img_array[18][13][13] <= img[8275];\
        in_img_array[18][13][14] <= img[8276];\
        in_img_array[18][13][15] <= img[8277];\
        in_img_array[18][13][16] <= img[8278];\
        in_img_array[18][13][17] <= img[8279];\
        in_img_array[18][14][0] <= img[8280];\
        in_img_array[18][14][1] <= img[8281];\
        in_img_array[18][14][2] <= img[8282];\
        in_img_array[18][14][3] <= img[8283];\
        in_img_array[18][14][4] <= img[8284];\
        in_img_array[18][14][5] <= img[8285];\
        in_img_array[18][14][6] <= img[8286];\
        in_img_array[18][14][7] <= img[8287];\
        in_img_array[18][14][8] <= img[8288];\
        in_img_array[18][14][9] <= img[8289];\
        in_img_array[18][14][10] <= img[8290];\
        in_img_array[18][14][11] <= img[8291];\
        in_img_array[18][14][12] <= img[8292];\
        in_img_array[18][14][13] <= img[8293];\
        in_img_array[18][14][14] <= img[8294];\
        in_img_array[18][14][15] <= img[8295];\
        in_img_array[18][14][16] <= img[8296];\
        in_img_array[18][14][17] <= img[8297];\
        in_img_array[18][15][0] <= img[8298];\
        in_img_array[18][15][1] <= img[8299];\
        in_img_array[18][15][2] <= img[8300];\
        in_img_array[18][15][3] <= img[8301];\
        in_img_array[18][15][4] <= img[8302];\
        in_img_array[18][15][5] <= img[8303];\
        in_img_array[18][15][6] <= img[8304];\
        in_img_array[18][15][7] <= img[8305];\
        in_img_array[18][15][8] <= img[8306];\
        in_img_array[18][15][9] <= img[8307];\
        in_img_array[18][15][10] <= img[8308];\
        in_img_array[18][15][11] <= img[8309];\
        in_img_array[18][15][12] <= img[8310];\
        in_img_array[18][15][13] <= img[8311];\
        in_img_array[18][15][14] <= img[8312];\
        in_img_array[18][15][15] <= img[8313];\
        in_img_array[18][15][16] <= img[8314];\
        in_img_array[18][15][17] <= img[8315];\
        in_img_array[18][16][0] <= img[8316];\
        in_img_array[18][16][1] <= img[8317];\
        in_img_array[18][16][2] <= img[8318];\
        in_img_array[18][16][3] <= img[8319];\
        in_img_array[18][16][4] <= img[8320];\
        in_img_array[18][16][5] <= img[8321];\
        in_img_array[18][16][6] <= img[8322];\
        in_img_array[18][16][7] <= img[8323];\
        in_img_array[18][16][8] <= img[8324];\
        in_img_array[18][16][9] <= img[8325];\
        in_img_array[18][16][10] <= img[8326];\
        in_img_array[18][16][11] <= img[8327];\
        in_img_array[18][16][12] <= img[8328];\
        in_img_array[18][16][13] <= img[8329];\
        in_img_array[18][16][14] <= img[8330];\
        in_img_array[18][16][15] <= img[8331];\
        in_img_array[18][16][16] <= img[8332];\
        in_img_array[18][16][17] <= img[8333];\
        in_img_array[18][17][0] <= img[8334];\
        in_img_array[18][17][1] <= img[8335];\
        in_img_array[18][17][2] <= img[8336];\
        in_img_array[18][17][3] <= img[8337];\
        in_img_array[18][17][4] <= img[8338];\
        in_img_array[18][17][5] <= img[8339];\
        in_img_array[18][17][6] <= img[8340];\
        in_img_array[18][17][7] <= img[8341];\
        in_img_array[18][17][8] <= img[8342];\
        in_img_array[18][17][9] <= img[8343];\
        in_img_array[18][17][10] <= img[8344];\
        in_img_array[18][17][11] <= img[8345];\
        in_img_array[18][17][12] <= img[8346];\
        in_img_array[18][17][13] <= img[8347];\
        in_img_array[18][17][14] <= img[8348];\
        in_img_array[18][17][15] <= img[8349];\
        in_img_array[18][17][16] <= img[8350];\
        in_img_array[18][17][17] <= img[8351];\
        in_img_array[18][18][0] <= img[8352];\
        in_img_array[18][18][1] <= img[8353];\
        in_img_array[18][18][2] <= img[8354];\
        in_img_array[18][18][3] <= img[8355];\
        in_img_array[18][18][4] <= img[8356];\
        in_img_array[18][18][5] <= img[8357];\
        in_img_array[18][18][6] <= img[8358];\
        in_img_array[18][18][7] <= img[8359];\
        in_img_array[18][18][8] <= img[8360];\
        in_img_array[18][18][9] <= img[8361];\
        in_img_array[18][18][10] <= img[8362];\
        in_img_array[18][18][11] <= img[8363];\
        in_img_array[18][18][12] <= img[8364];\
        in_img_array[18][18][13] <= img[8365];\
        in_img_array[18][18][14] <= img[8366];\
        in_img_array[18][18][15] <= img[8367];\
        in_img_array[18][18][16] <= img[8368];\
        in_img_array[18][18][17] <= img[8369];\
        in_img_array[18][19][0] <= img[8370];\
        in_img_array[18][19][1] <= img[8371];\
        in_img_array[18][19][2] <= img[8372];\
        in_img_array[18][19][3] <= img[8373];\
        in_img_array[18][19][4] <= img[8374];\
        in_img_array[18][19][5] <= img[8375];\
        in_img_array[18][19][6] <= img[8376];\
        in_img_array[18][19][7] <= img[8377];\
        in_img_array[18][19][8] <= img[8378];\
        in_img_array[18][19][9] <= img[8379];\
        in_img_array[18][19][10] <= img[8380];\
        in_img_array[18][19][11] <= img[8381];\
        in_img_array[18][19][12] <= img[8382];\
        in_img_array[18][19][13] <= img[8383];\
        in_img_array[18][19][14] <= img[8384];\
        in_img_array[18][19][15] <= img[8385];\
        in_img_array[18][19][16] <= img[8386];\
        in_img_array[18][19][17] <= img[8387];\
        in_img_array[18][20][0] <= img[8388];\
        in_img_array[18][20][1] <= img[8389];\
        in_img_array[18][20][2] <= img[8390];\
        in_img_array[18][20][3] <= img[8391];\
        in_img_array[18][20][4] <= img[8392];\
        in_img_array[18][20][5] <= img[8393];\
        in_img_array[18][20][6] <= img[8394];\
        in_img_array[18][20][7] <= img[8395];\
        in_img_array[18][20][8] <= img[8396];\
        in_img_array[18][20][9] <= img[8397];\
        in_img_array[18][20][10] <= img[8398];\
        in_img_array[18][20][11] <= img[8399];\
        in_img_array[18][20][12] <= img[8400];\
        in_img_array[18][20][13] <= img[8401];\
        in_img_array[18][20][14] <= img[8402];\
        in_img_array[18][20][15] <= img[8403];\
        in_img_array[18][20][16] <= img[8404];\
        in_img_array[18][20][17] <= img[8405];\
        in_img_array[18][21][0] <= img[8406];\
        in_img_array[18][21][1] <= img[8407];\
        in_img_array[18][21][2] <= img[8408];\
        in_img_array[18][21][3] <= img[8409];\
        in_img_array[18][21][4] <= img[8410];\
        in_img_array[18][21][5] <= img[8411];\
        in_img_array[18][21][6] <= img[8412];\
        in_img_array[18][21][7] <= img[8413];\
        in_img_array[18][21][8] <= img[8414];\
        in_img_array[18][21][9] <= img[8415];\
        in_img_array[18][21][10] <= img[8416];\
        in_img_array[18][21][11] <= img[8417];\
        in_img_array[18][21][12] <= img[8418];\
        in_img_array[18][21][13] <= img[8419];\
        in_img_array[18][21][14] <= img[8420];\
        in_img_array[18][21][15] <= img[8421];\
        in_img_array[18][21][16] <= img[8422];\
        in_img_array[18][21][17] <= img[8423];\
        in_img_array[18][22][0] <= img[8424];\
        in_img_array[18][22][1] <= img[8425];\
        in_img_array[18][22][2] <= img[8426];\
        in_img_array[18][22][3] <= img[8427];\
        in_img_array[18][22][4] <= img[8428];\
        in_img_array[18][22][5] <= img[8429];\
        in_img_array[18][22][6] <= img[8430];\
        in_img_array[18][22][7] <= img[8431];\
        in_img_array[18][22][8] <= img[8432];\
        in_img_array[18][22][9] <= img[8433];\
        in_img_array[18][22][10] <= img[8434];\
        in_img_array[18][22][11] <= img[8435];\
        in_img_array[18][22][12] <= img[8436];\
        in_img_array[18][22][13] <= img[8437];\
        in_img_array[18][22][14] <= img[8438];\
        in_img_array[18][22][15] <= img[8439];\
        in_img_array[18][22][16] <= img[8440];\
        in_img_array[18][22][17] <= img[8441];\
        in_img_array[18][23][0] <= img[8442];\
        in_img_array[18][23][1] <= img[8443];\
        in_img_array[18][23][2] <= img[8444];\
        in_img_array[18][23][3] <= img[8445];\
        in_img_array[18][23][4] <= img[8446];\
        in_img_array[18][23][5] <= img[8447];\
        in_img_array[18][23][6] <= img[8448];\
        in_img_array[18][23][7] <= img[8449];\
        in_img_array[18][23][8] <= img[8450];\
        in_img_array[18][23][9] <= img[8451];\
        in_img_array[18][23][10] <= img[8452];\
        in_img_array[18][23][11] <= img[8453];\
        in_img_array[18][23][12] <= img[8454];\
        in_img_array[18][23][13] <= img[8455];\
        in_img_array[18][23][14] <= img[8456];\
        in_img_array[18][23][15] <= img[8457];\
        in_img_array[18][23][16] <= img[8458];\
        in_img_array[18][23][17] <= img[8459];\
        in_img_array[18][24][0] <= img[8460];\
        in_img_array[18][24][1] <= img[8461];\
        in_img_array[18][24][2] <= img[8462];\
        in_img_array[18][24][3] <= img[8463];\
        in_img_array[18][24][4] <= img[8464];\
        in_img_array[18][24][5] <= img[8465];\
        in_img_array[18][24][6] <= img[8466];\
        in_img_array[18][24][7] <= img[8467];\
        in_img_array[18][24][8] <= img[8468];\
        in_img_array[18][24][9] <= img[8469];\
        in_img_array[18][24][10] <= img[8470];\
        in_img_array[18][24][11] <= img[8471];\
        in_img_array[18][24][12] <= img[8472];\
        in_img_array[18][24][13] <= img[8473];\
        in_img_array[18][24][14] <= img[8474];\
        in_img_array[18][24][15] <= img[8475];\
        in_img_array[18][24][16] <= img[8476];\
        in_img_array[18][24][17] <= img[8477];\
        in_img_array[18][25][0] <= img[8478];\
        in_img_array[18][25][1] <= img[8479];\
        in_img_array[18][25][2] <= img[8480];\
        in_img_array[18][25][3] <= img[8481];\
        in_img_array[18][25][4] <= img[8482];\
        in_img_array[18][25][5] <= img[8483];\
        in_img_array[18][25][6] <= img[8484];\
        in_img_array[18][25][7] <= img[8485];\
        in_img_array[18][25][8] <= img[8486];\
        in_img_array[18][25][9] <= img[8487];\
        in_img_array[18][25][10] <= img[8488];\
        in_img_array[18][25][11] <= img[8489];\
        in_img_array[18][25][12] <= img[8490];\
        in_img_array[18][25][13] <= img[8491];\
        in_img_array[18][25][14] <= img[8492];\
        in_img_array[18][25][15] <= img[8493];\
        in_img_array[18][25][16] <= img[8494];\
        in_img_array[18][25][17] <= img[8495];\
        in_img_array[18][26][0] <= img[8496];\
        in_img_array[18][26][1] <= img[8497];\
        in_img_array[18][26][2] <= img[8498];\
        in_img_array[18][26][3] <= img[8499];\
        in_img_array[18][26][4] <= img[8500];\
        in_img_array[18][26][5] <= img[8501];\
        in_img_array[18][26][6] <= img[8502];\
        in_img_array[18][26][7] <= img[8503];\
        in_img_array[18][26][8] <= img[8504];\
        in_img_array[18][26][9] <= img[8505];\
        in_img_array[18][26][10] <= img[8506];\
        in_img_array[18][26][11] <= img[8507];\
        in_img_array[18][26][12] <= img[8508];\
        in_img_array[18][26][13] <= img[8509];\
        in_img_array[18][26][14] <= img[8510];\
        in_img_array[18][26][15] <= img[8511];\
        in_img_array[18][26][16] <= img[8512];\
        in_img_array[18][26][17] <= img[8513];\
        in_img_array[18][27][0] <= img[8514];\
        in_img_array[18][27][1] <= img[8515];\
        in_img_array[18][27][2] <= img[8516];\
        in_img_array[18][27][3] <= img[8517];\
        in_img_array[18][27][4] <= img[8518];\
        in_img_array[18][27][5] <= img[8519];\
        in_img_array[18][27][6] <= img[8520];\
        in_img_array[18][27][7] <= img[8521];\
        in_img_array[18][27][8] <= img[8522];\
        in_img_array[18][27][9] <= img[8523];\
        in_img_array[18][27][10] <= img[8524];\
        in_img_array[18][27][11] <= img[8525];\
        in_img_array[18][27][12] <= img[8526];\
        in_img_array[18][27][13] <= img[8527];\
        in_img_array[18][27][14] <= img[8528];\
        in_img_array[18][27][15] <= img[8529];\
        in_img_array[18][27][16] <= img[8530];\
        in_img_array[18][27][17] <= img[8531];\
        in_img_array[18][28][0] <= img[8532];\
        in_img_array[18][28][1] <= img[8533];\
        in_img_array[18][28][2] <= img[8534];\
        in_img_array[18][28][3] <= img[8535];\
        in_img_array[18][28][4] <= img[8536];\
        in_img_array[18][28][5] <= img[8537];\
        in_img_array[18][28][6] <= img[8538];\
        in_img_array[18][28][7] <= img[8539];\
        in_img_array[18][28][8] <= img[8540];\
        in_img_array[18][28][9] <= img[8541];\
        in_img_array[18][28][10] <= img[8542];\
        in_img_array[18][28][11] <= img[8543];\
        in_img_array[18][28][12] <= img[8544];\
        in_img_array[18][28][13] <= img[8545];\
        in_img_array[18][28][14] <= img[8546];\
        in_img_array[18][28][15] <= img[8547];\
        in_img_array[18][28][16] <= img[8548];\
        in_img_array[18][28][17] <= img[8549];\
        in_img_array[18][29][0] <= img[8550];\
        in_img_array[18][29][1] <= img[8551];\
        in_img_array[18][29][2] <= img[8552];\
        in_img_array[18][29][3] <= img[8553];\
        in_img_array[18][29][4] <= img[8554];\
        in_img_array[18][29][5] <= img[8555];\
        in_img_array[18][29][6] <= img[8556];\
        in_img_array[18][29][7] <= img[8557];\
        in_img_array[18][29][8] <= img[8558];\
        in_img_array[18][29][9] <= img[8559];\
        in_img_array[18][29][10] <= img[8560];\
        in_img_array[18][29][11] <= img[8561];\
        in_img_array[18][29][12] <= img[8562];\
        in_img_array[18][29][13] <= img[8563];\
        in_img_array[18][29][14] <= img[8564];\
        in_img_array[18][29][15] <= img[8565];\
        in_img_array[18][29][16] <= img[8566];\
        in_img_array[18][29][17] <= img[8567];\
        in_img_array[19][2][0] <= img[8568];\
        in_img_array[19][2][1] <= img[8569];\
        in_img_array[19][2][2] <= img[8570];\
        in_img_array[19][2][3] <= img[8571];\
        in_img_array[19][2][4] <= img[8572];\
        in_img_array[19][2][5] <= img[8573];\
        in_img_array[19][2][6] <= img[8574];\
        in_img_array[19][2][7] <= img[8575];\
        in_img_array[19][2][8] <= img[8576];\
        in_img_array[19][2][9] <= img[8577];\
        in_img_array[19][2][10] <= img[8578];\
        in_img_array[19][2][11] <= img[8579];\
        in_img_array[19][2][12] <= img[8580];\
        in_img_array[19][2][13] <= img[8581];\
        in_img_array[19][2][14] <= img[8582];\
        in_img_array[19][2][15] <= img[8583];\
        in_img_array[19][2][16] <= img[8584];\
        in_img_array[19][2][17] <= img[8585];\
        in_img_array[19][3][0] <= img[8586];\
        in_img_array[19][3][1] <= img[8587];\
        in_img_array[19][3][2] <= img[8588];\
        in_img_array[19][3][3] <= img[8589];\
        in_img_array[19][3][4] <= img[8590];\
        in_img_array[19][3][5] <= img[8591];\
        in_img_array[19][3][6] <= img[8592];\
        in_img_array[19][3][7] <= img[8593];\
        in_img_array[19][3][8] <= img[8594];\
        in_img_array[19][3][9] <= img[8595];\
        in_img_array[19][3][10] <= img[8596];\
        in_img_array[19][3][11] <= img[8597];\
        in_img_array[19][3][12] <= img[8598];\
        in_img_array[19][3][13] <= img[8599];\
        in_img_array[19][3][14] <= img[8600];\
        in_img_array[19][3][15] <= img[8601];\
        in_img_array[19][3][16] <= img[8602];\
        in_img_array[19][3][17] <= img[8603];\
        in_img_array[19][4][0] <= img[8604];\
        in_img_array[19][4][1] <= img[8605];\
        in_img_array[19][4][2] <= img[8606];\
        in_img_array[19][4][3] <= img[8607];\
        in_img_array[19][4][4] <= img[8608];\
        in_img_array[19][4][5] <= img[8609];\
        in_img_array[19][4][6] <= img[8610];\
        in_img_array[19][4][7] <= img[8611];\
        in_img_array[19][4][8] <= img[8612];\
        in_img_array[19][4][9] <= img[8613];\
        in_img_array[19][4][10] <= img[8614];\
        in_img_array[19][4][11] <= img[8615];\
        in_img_array[19][4][12] <= img[8616];\
        in_img_array[19][4][13] <= img[8617];\
        in_img_array[19][4][14] <= img[8618];\
        in_img_array[19][4][15] <= img[8619];\
        in_img_array[19][4][16] <= img[8620];\
        in_img_array[19][4][17] <= img[8621];\
        in_img_array[19][5][0] <= img[8622];\
        in_img_array[19][5][1] <= img[8623];\
        in_img_array[19][5][2] <= img[8624];\
        in_img_array[19][5][3] <= img[8625];\
        in_img_array[19][5][4] <= img[8626];\
        in_img_array[19][5][5] <= img[8627];\
        in_img_array[19][5][6] <= img[8628];\
        in_img_array[19][5][7] <= img[8629];\
        in_img_array[19][5][8] <= img[8630];\
        in_img_array[19][5][9] <= img[8631];\
        in_img_array[19][5][10] <= img[8632];\
        in_img_array[19][5][11] <= img[8633];\
        in_img_array[19][5][12] <= img[8634];\
        in_img_array[19][5][13] <= img[8635];\
        in_img_array[19][5][14] <= img[8636];\
        in_img_array[19][5][15] <= img[8637];\
        in_img_array[19][5][16] <= img[8638];\
        in_img_array[19][5][17] <= img[8639];\
        in_img_array[19][6][0] <= img[8640];\
        in_img_array[19][6][1] <= img[8641];\
        in_img_array[19][6][2] <= img[8642];\
        in_img_array[19][6][3] <= img[8643];\
        in_img_array[19][6][4] <= img[8644];\
        in_img_array[19][6][5] <= img[8645];\
        in_img_array[19][6][6] <= img[8646];\
        in_img_array[19][6][7] <= img[8647];\
        in_img_array[19][6][8] <= img[8648];\
        in_img_array[19][6][9] <= img[8649];\
        in_img_array[19][6][10] <= img[8650];\
        in_img_array[19][6][11] <= img[8651];\
        in_img_array[19][6][12] <= img[8652];\
        in_img_array[19][6][13] <= img[8653];\
        in_img_array[19][6][14] <= img[8654];\
        in_img_array[19][6][15] <= img[8655];\
        in_img_array[19][6][16] <= img[8656];\
        in_img_array[19][6][17] <= img[8657];\
        in_img_array[19][7][0] <= img[8658];\
        in_img_array[19][7][1] <= img[8659];\
        in_img_array[19][7][2] <= img[8660];\
        in_img_array[19][7][3] <= img[8661];\
        in_img_array[19][7][4] <= img[8662];\
        in_img_array[19][7][5] <= img[8663];\
        in_img_array[19][7][6] <= img[8664];\
        in_img_array[19][7][7] <= img[8665];\
        in_img_array[19][7][8] <= img[8666];\
        in_img_array[19][7][9] <= img[8667];\
        in_img_array[19][7][10] <= img[8668];\
        in_img_array[19][7][11] <= img[8669];\
        in_img_array[19][7][12] <= img[8670];\
        in_img_array[19][7][13] <= img[8671];\
        in_img_array[19][7][14] <= img[8672];\
        in_img_array[19][7][15] <= img[8673];\
        in_img_array[19][7][16] <= img[8674];\
        in_img_array[19][7][17] <= img[8675];\
        in_img_array[19][8][0] <= img[8676];\
        in_img_array[19][8][1] <= img[8677];\
        in_img_array[19][8][2] <= img[8678];\
        in_img_array[19][8][3] <= img[8679];\
        in_img_array[19][8][4] <= img[8680];\
        in_img_array[19][8][5] <= img[8681];\
        in_img_array[19][8][6] <= img[8682];\
        in_img_array[19][8][7] <= img[8683];\
        in_img_array[19][8][8] <= img[8684];\
        in_img_array[19][8][9] <= img[8685];\
        in_img_array[19][8][10] <= img[8686];\
        in_img_array[19][8][11] <= img[8687];\
        in_img_array[19][8][12] <= img[8688];\
        in_img_array[19][8][13] <= img[8689];\
        in_img_array[19][8][14] <= img[8690];\
        in_img_array[19][8][15] <= img[8691];\
        in_img_array[19][8][16] <= img[8692];\
        in_img_array[19][8][17] <= img[8693];\
        in_img_array[19][9][0] <= img[8694];\
        in_img_array[19][9][1] <= img[8695];\
        in_img_array[19][9][2] <= img[8696];\
        in_img_array[19][9][3] <= img[8697];\
        in_img_array[19][9][4] <= img[8698];\
        in_img_array[19][9][5] <= img[8699];\
        in_img_array[19][9][6] <= img[8700];\
        in_img_array[19][9][7] <= img[8701];\
        in_img_array[19][9][8] <= img[8702];\
        in_img_array[19][9][9] <= img[8703];\
        in_img_array[19][9][10] <= img[8704];\
        in_img_array[19][9][11] <= img[8705];\
        in_img_array[19][9][12] <= img[8706];\
        in_img_array[19][9][13] <= img[8707];\
        in_img_array[19][9][14] <= img[8708];\
        in_img_array[19][9][15] <= img[8709];\
        in_img_array[19][9][16] <= img[8710];\
        in_img_array[19][9][17] <= img[8711];\
        in_img_array[19][10][0] <= img[8712];\
        in_img_array[19][10][1] <= img[8713];\
        in_img_array[19][10][2] <= img[8714];\
        in_img_array[19][10][3] <= img[8715];\
        in_img_array[19][10][4] <= img[8716];\
        in_img_array[19][10][5] <= img[8717];\
        in_img_array[19][10][6] <= img[8718];\
        in_img_array[19][10][7] <= img[8719];\
        in_img_array[19][10][8] <= img[8720];\
        in_img_array[19][10][9] <= img[8721];\
        in_img_array[19][10][10] <= img[8722];\
        in_img_array[19][10][11] <= img[8723];\
        in_img_array[19][10][12] <= img[8724];\
        in_img_array[19][10][13] <= img[8725];\
        in_img_array[19][10][14] <= img[8726];\
        in_img_array[19][10][15] <= img[8727];\
        in_img_array[19][10][16] <= img[8728];\
        in_img_array[19][10][17] <= img[8729];\
        in_img_array[19][11][0] <= img[8730];\
        in_img_array[19][11][1] <= img[8731];\
        in_img_array[19][11][2] <= img[8732];\
        in_img_array[19][11][3] <= img[8733];\
        in_img_array[19][11][4] <= img[8734];\
        in_img_array[19][11][5] <= img[8735];\
        in_img_array[19][11][6] <= img[8736];\
        in_img_array[19][11][7] <= img[8737];\
        in_img_array[19][11][8] <= img[8738];\
        in_img_array[19][11][9] <= img[8739];\
        in_img_array[19][11][10] <= img[8740];\
        in_img_array[19][11][11] <= img[8741];\
        in_img_array[19][11][12] <= img[8742];\
        in_img_array[19][11][13] <= img[8743];\
        in_img_array[19][11][14] <= img[8744];\
        in_img_array[19][11][15] <= img[8745];\
        in_img_array[19][11][16] <= img[8746];\
        in_img_array[19][11][17] <= img[8747];\
        in_img_array[19][12][0] <= img[8748];\
        in_img_array[19][12][1] <= img[8749];\
        in_img_array[19][12][2] <= img[8750];\
        in_img_array[19][12][3] <= img[8751];\
        in_img_array[19][12][4] <= img[8752];\
        in_img_array[19][12][5] <= img[8753];\
        in_img_array[19][12][6] <= img[8754];\
        in_img_array[19][12][7] <= img[8755];\
        in_img_array[19][12][8] <= img[8756];\
        in_img_array[19][12][9] <= img[8757];\
        in_img_array[19][12][10] <= img[8758];\
        in_img_array[19][12][11] <= img[8759];\
        in_img_array[19][12][12] <= img[8760];\
        in_img_array[19][12][13] <= img[8761];\
        in_img_array[19][12][14] <= img[8762];\
        in_img_array[19][12][15] <= img[8763];\
        in_img_array[19][12][16] <= img[8764];\
        in_img_array[19][12][17] <= img[8765];\
        in_img_array[19][13][0] <= img[8766];\
        in_img_array[19][13][1] <= img[8767];\
        in_img_array[19][13][2] <= img[8768];\
        in_img_array[19][13][3] <= img[8769];\
        in_img_array[19][13][4] <= img[8770];\
        in_img_array[19][13][5] <= img[8771];\
        in_img_array[19][13][6] <= img[8772];\
        in_img_array[19][13][7] <= img[8773];\
        in_img_array[19][13][8] <= img[8774];\
        in_img_array[19][13][9] <= img[8775];\
        in_img_array[19][13][10] <= img[8776];\
        in_img_array[19][13][11] <= img[8777];\
        in_img_array[19][13][12] <= img[8778];\
        in_img_array[19][13][13] <= img[8779];\
        in_img_array[19][13][14] <= img[8780];\
        in_img_array[19][13][15] <= img[8781];\
        in_img_array[19][13][16] <= img[8782];\
        in_img_array[19][13][17] <= img[8783];\
        in_img_array[19][14][0] <= img[8784];\
        in_img_array[19][14][1] <= img[8785];\
        in_img_array[19][14][2] <= img[8786];\
        in_img_array[19][14][3] <= img[8787];\
        in_img_array[19][14][4] <= img[8788];\
        in_img_array[19][14][5] <= img[8789];\
        in_img_array[19][14][6] <= img[8790];\
        in_img_array[19][14][7] <= img[8791];\
        in_img_array[19][14][8] <= img[8792];\
        in_img_array[19][14][9] <= img[8793];\
        in_img_array[19][14][10] <= img[8794];\
        in_img_array[19][14][11] <= img[8795];\
        in_img_array[19][14][12] <= img[8796];\
        in_img_array[19][14][13] <= img[8797];\
        in_img_array[19][14][14] <= img[8798];\
        in_img_array[19][14][15] <= img[8799];\
        in_img_array[19][14][16] <= img[8800];\
        in_img_array[19][14][17] <= img[8801];\
        in_img_array[19][15][0] <= img[8802];\
        in_img_array[19][15][1] <= img[8803];\
        in_img_array[19][15][2] <= img[8804];\
        in_img_array[19][15][3] <= img[8805];\
        in_img_array[19][15][4] <= img[8806];\
        in_img_array[19][15][5] <= img[8807];\
        in_img_array[19][15][6] <= img[8808];\
        in_img_array[19][15][7] <= img[8809];\
        in_img_array[19][15][8] <= img[8810];\
        in_img_array[19][15][9] <= img[8811];\
        in_img_array[19][15][10] <= img[8812];\
        in_img_array[19][15][11] <= img[8813];\
        in_img_array[19][15][12] <= img[8814];\
        in_img_array[19][15][13] <= img[8815];\
        in_img_array[19][15][14] <= img[8816];\
        in_img_array[19][15][15] <= img[8817];\
        in_img_array[19][15][16] <= img[8818];\
        in_img_array[19][15][17] <= img[8819];\
        in_img_array[19][16][0] <= img[8820];\
        in_img_array[19][16][1] <= img[8821];\
        in_img_array[19][16][2] <= img[8822];\
        in_img_array[19][16][3] <= img[8823];\
        in_img_array[19][16][4] <= img[8824];\
        in_img_array[19][16][5] <= img[8825];\
        in_img_array[19][16][6] <= img[8826];\
        in_img_array[19][16][7] <= img[8827];\
        in_img_array[19][16][8] <= img[8828];\
        in_img_array[19][16][9] <= img[8829];\
        in_img_array[19][16][10] <= img[8830];\
        in_img_array[19][16][11] <= img[8831];\
        in_img_array[19][16][12] <= img[8832];\
        in_img_array[19][16][13] <= img[8833];\
        in_img_array[19][16][14] <= img[8834];\
        in_img_array[19][16][15] <= img[8835];\
        in_img_array[19][16][16] <= img[8836];\
        in_img_array[19][16][17] <= img[8837];\
        in_img_array[19][17][0] <= img[8838];\
        in_img_array[19][17][1] <= img[8839];\
        in_img_array[19][17][2] <= img[8840];\
        in_img_array[19][17][3] <= img[8841];\
        in_img_array[19][17][4] <= img[8842];\
        in_img_array[19][17][5] <= img[8843];\
        in_img_array[19][17][6] <= img[8844];\
        in_img_array[19][17][7] <= img[8845];\
        in_img_array[19][17][8] <= img[8846];\
        in_img_array[19][17][9] <= img[8847];\
        in_img_array[19][17][10] <= img[8848];\
        in_img_array[19][17][11] <= img[8849];\
        in_img_array[19][17][12] <= img[8850];\
        in_img_array[19][17][13] <= img[8851];\
        in_img_array[19][17][14] <= img[8852];\
        in_img_array[19][17][15] <= img[8853];\
        in_img_array[19][17][16] <= img[8854];\
        in_img_array[19][17][17] <= img[8855];\
        in_img_array[19][18][0] <= img[8856];\
        in_img_array[19][18][1] <= img[8857];\
        in_img_array[19][18][2] <= img[8858];\
        in_img_array[19][18][3] <= img[8859];\
        in_img_array[19][18][4] <= img[8860];\
        in_img_array[19][18][5] <= img[8861];\
        in_img_array[19][18][6] <= img[8862];\
        in_img_array[19][18][7] <= img[8863];\
        in_img_array[19][18][8] <= img[8864];\
        in_img_array[19][18][9] <= img[8865];\
        in_img_array[19][18][10] <= img[8866];\
        in_img_array[19][18][11] <= img[8867];\
        in_img_array[19][18][12] <= img[8868];\
        in_img_array[19][18][13] <= img[8869];\
        in_img_array[19][18][14] <= img[8870];\
        in_img_array[19][18][15] <= img[8871];\
        in_img_array[19][18][16] <= img[8872];\
        in_img_array[19][18][17] <= img[8873];\
        in_img_array[19][19][0] <= img[8874];\
        in_img_array[19][19][1] <= img[8875];\
        in_img_array[19][19][2] <= img[8876];\
        in_img_array[19][19][3] <= img[8877];\
        in_img_array[19][19][4] <= img[8878];\
        in_img_array[19][19][5] <= img[8879];\
        in_img_array[19][19][6] <= img[8880];\
        in_img_array[19][19][7] <= img[8881];\
        in_img_array[19][19][8] <= img[8882];\
        in_img_array[19][19][9] <= img[8883];\
        in_img_array[19][19][10] <= img[8884];\
        in_img_array[19][19][11] <= img[8885];\
        in_img_array[19][19][12] <= img[8886];\
        in_img_array[19][19][13] <= img[8887];\
        in_img_array[19][19][14] <= img[8888];\
        in_img_array[19][19][15] <= img[8889];\
        in_img_array[19][19][16] <= img[8890];\
        in_img_array[19][19][17] <= img[8891];\
        in_img_array[19][20][0] <= img[8892];\
        in_img_array[19][20][1] <= img[8893];\
        in_img_array[19][20][2] <= img[8894];\
        in_img_array[19][20][3] <= img[8895];\
        in_img_array[19][20][4] <= img[8896];\
        in_img_array[19][20][5] <= img[8897];\
        in_img_array[19][20][6] <= img[8898];\
        in_img_array[19][20][7] <= img[8899];\
        in_img_array[19][20][8] <= img[8900];\
        in_img_array[19][20][9] <= img[8901];\
        in_img_array[19][20][10] <= img[8902];\
        in_img_array[19][20][11] <= img[8903];\
        in_img_array[19][20][12] <= img[8904];\
        in_img_array[19][20][13] <= img[8905];\
        in_img_array[19][20][14] <= img[8906];\
        in_img_array[19][20][15] <= img[8907];\
        in_img_array[19][20][16] <= img[8908];\
        in_img_array[19][20][17] <= img[8909];\
        in_img_array[19][21][0] <= img[8910];\
        in_img_array[19][21][1] <= img[8911];\
        in_img_array[19][21][2] <= img[8912];\
        in_img_array[19][21][3] <= img[8913];\
        in_img_array[19][21][4] <= img[8914];\
        in_img_array[19][21][5] <= img[8915];\
        in_img_array[19][21][6] <= img[8916];\
        in_img_array[19][21][7] <= img[8917];\
        in_img_array[19][21][8] <= img[8918];\
        in_img_array[19][21][9] <= img[8919];\
        in_img_array[19][21][10] <= img[8920];\
        in_img_array[19][21][11] <= img[8921];\
        in_img_array[19][21][12] <= img[8922];\
        in_img_array[19][21][13] <= img[8923];\
        in_img_array[19][21][14] <= img[8924];\
        in_img_array[19][21][15] <= img[8925];\
        in_img_array[19][21][16] <= img[8926];\
        in_img_array[19][21][17] <= img[8927];\
        in_img_array[19][22][0] <= img[8928];\
        in_img_array[19][22][1] <= img[8929];\
        in_img_array[19][22][2] <= img[8930];\
        in_img_array[19][22][3] <= img[8931];\
        in_img_array[19][22][4] <= img[8932];\
        in_img_array[19][22][5] <= img[8933];\
        in_img_array[19][22][6] <= img[8934];\
        in_img_array[19][22][7] <= img[8935];\
        in_img_array[19][22][8] <= img[8936];\
        in_img_array[19][22][9] <= img[8937];\
        in_img_array[19][22][10] <= img[8938];\
        in_img_array[19][22][11] <= img[8939];\
        in_img_array[19][22][12] <= img[8940];\
        in_img_array[19][22][13] <= img[8941];\
        in_img_array[19][22][14] <= img[8942];\
        in_img_array[19][22][15] <= img[8943];\
        in_img_array[19][22][16] <= img[8944];\
        in_img_array[19][22][17] <= img[8945];\
        in_img_array[19][23][0] <= img[8946];\
        in_img_array[19][23][1] <= img[8947];\
        in_img_array[19][23][2] <= img[8948];\
        in_img_array[19][23][3] <= img[8949];\
        in_img_array[19][23][4] <= img[8950];\
        in_img_array[19][23][5] <= img[8951];\
        in_img_array[19][23][6] <= img[8952];\
        in_img_array[19][23][7] <= img[8953];\
        in_img_array[19][23][8] <= img[8954];\
        in_img_array[19][23][9] <= img[8955];\
        in_img_array[19][23][10] <= img[8956];\
        in_img_array[19][23][11] <= img[8957];\
        in_img_array[19][23][12] <= img[8958];\
        in_img_array[19][23][13] <= img[8959];\
        in_img_array[19][23][14] <= img[8960];\
        in_img_array[19][23][15] <= img[8961];\
        in_img_array[19][23][16] <= img[8962];\
        in_img_array[19][23][17] <= img[8963];\
        in_img_array[19][24][0] <= img[8964];\
        in_img_array[19][24][1] <= img[8965];\
        in_img_array[19][24][2] <= img[8966];\
        in_img_array[19][24][3] <= img[8967];\
        in_img_array[19][24][4] <= img[8968];\
        in_img_array[19][24][5] <= img[8969];\
        in_img_array[19][24][6] <= img[8970];\
        in_img_array[19][24][7] <= img[8971];\
        in_img_array[19][24][8] <= img[8972];\
        in_img_array[19][24][9] <= img[8973];\
        in_img_array[19][24][10] <= img[8974];\
        in_img_array[19][24][11] <= img[8975];\
        in_img_array[19][24][12] <= img[8976];\
        in_img_array[19][24][13] <= img[8977];\
        in_img_array[19][24][14] <= img[8978];\
        in_img_array[19][24][15] <= img[8979];\
        in_img_array[19][24][16] <= img[8980];\
        in_img_array[19][24][17] <= img[8981];\
        in_img_array[19][25][0] <= img[8982];\
        in_img_array[19][25][1] <= img[8983];\
        in_img_array[19][25][2] <= img[8984];\
        in_img_array[19][25][3] <= img[8985];\
        in_img_array[19][25][4] <= img[8986];\
        in_img_array[19][25][5] <= img[8987];\
        in_img_array[19][25][6] <= img[8988];\
        in_img_array[19][25][7] <= img[8989];\
        in_img_array[19][25][8] <= img[8990];\
        in_img_array[19][25][9] <= img[8991];\
        in_img_array[19][25][10] <= img[8992];\
        in_img_array[19][25][11] <= img[8993];\
        in_img_array[19][25][12] <= img[8994];\
        in_img_array[19][25][13] <= img[8995];\
        in_img_array[19][25][14] <= img[8996];\
        in_img_array[19][25][15] <= img[8997];\
        in_img_array[19][25][16] <= img[8998];\
        in_img_array[19][25][17] <= img[8999];\
        in_img_array[19][26][0] <= img[9000];\
        in_img_array[19][26][1] <= img[9001];\
        in_img_array[19][26][2] <= img[9002];\
        in_img_array[19][26][3] <= img[9003];\
        in_img_array[19][26][4] <= img[9004];\
        in_img_array[19][26][5] <= img[9005];\
        in_img_array[19][26][6] <= img[9006];\
        in_img_array[19][26][7] <= img[9007];\
        in_img_array[19][26][8] <= img[9008];\
        in_img_array[19][26][9] <= img[9009];\
        in_img_array[19][26][10] <= img[9010];\
        in_img_array[19][26][11] <= img[9011];\
        in_img_array[19][26][12] <= img[9012];\
        in_img_array[19][26][13] <= img[9013];\
        in_img_array[19][26][14] <= img[9014];\
        in_img_array[19][26][15] <= img[9015];\
        in_img_array[19][26][16] <= img[9016];\
        in_img_array[19][26][17] <= img[9017];\
        in_img_array[19][27][0] <= img[9018];\
        in_img_array[19][27][1] <= img[9019];\
        in_img_array[19][27][2] <= img[9020];\
        in_img_array[19][27][3] <= img[9021];\
        in_img_array[19][27][4] <= img[9022];\
        in_img_array[19][27][5] <= img[9023];\
        in_img_array[19][27][6] <= img[9024];\
        in_img_array[19][27][7] <= img[9025];\
        in_img_array[19][27][8] <= img[9026];\
        in_img_array[19][27][9] <= img[9027];\
        in_img_array[19][27][10] <= img[9028];\
        in_img_array[19][27][11] <= img[9029];\
        in_img_array[19][27][12] <= img[9030];\
        in_img_array[19][27][13] <= img[9031];\
        in_img_array[19][27][14] <= img[9032];\
        in_img_array[19][27][15] <= img[9033];\
        in_img_array[19][27][16] <= img[9034];\
        in_img_array[19][27][17] <= img[9035];\
        in_img_array[19][28][0] <= img[9036];\
        in_img_array[19][28][1] <= img[9037];\
        in_img_array[19][28][2] <= img[9038];\
        in_img_array[19][28][3] <= img[9039];\
        in_img_array[19][28][4] <= img[9040];\
        in_img_array[19][28][5] <= img[9041];\
        in_img_array[19][28][6] <= img[9042];\
        in_img_array[19][28][7] <= img[9043];\
        in_img_array[19][28][8] <= img[9044];\
        in_img_array[19][28][9] <= img[9045];\
        in_img_array[19][28][10] <= img[9046];\
        in_img_array[19][28][11] <= img[9047];\
        in_img_array[19][28][12] <= img[9048];\
        in_img_array[19][28][13] <= img[9049];\
        in_img_array[19][28][14] <= img[9050];\
        in_img_array[19][28][15] <= img[9051];\
        in_img_array[19][28][16] <= img[9052];\
        in_img_array[19][28][17] <= img[9053];\
        in_img_array[19][29][0] <= img[9054];\
        in_img_array[19][29][1] <= img[9055];\
        in_img_array[19][29][2] <= img[9056];\
        in_img_array[19][29][3] <= img[9057];\
        in_img_array[19][29][4] <= img[9058];\
        in_img_array[19][29][5] <= img[9059];\
        in_img_array[19][29][6] <= img[9060];\
        in_img_array[19][29][7] <= img[9061];\
        in_img_array[19][29][8] <= img[9062];\
        in_img_array[19][29][9] <= img[9063];\
        in_img_array[19][29][10] <= img[9064];\
        in_img_array[19][29][11] <= img[9065];\
        in_img_array[19][29][12] <= img[9066];\
        in_img_array[19][29][13] <= img[9067];\
        in_img_array[19][29][14] <= img[9068];\
        in_img_array[19][29][15] <= img[9069];\
        in_img_array[19][29][16] <= img[9070];\
        in_img_array[19][29][17] <= img[9071];\
        in_img_array[20][2][0] <= img[9072];\
        in_img_array[20][2][1] <= img[9073];\
        in_img_array[20][2][2] <= img[9074];\
        in_img_array[20][2][3] <= img[9075];\
        in_img_array[20][2][4] <= img[9076];\
        in_img_array[20][2][5] <= img[9077];\
        in_img_array[20][2][6] <= img[9078];\
        in_img_array[20][2][7] <= img[9079];\
        in_img_array[20][2][8] <= img[9080];\
        in_img_array[20][2][9] <= img[9081];\
        in_img_array[20][2][10] <= img[9082];\
        in_img_array[20][2][11] <= img[9083];\
        in_img_array[20][2][12] <= img[9084];\
        in_img_array[20][2][13] <= img[9085];\
        in_img_array[20][2][14] <= img[9086];\
        in_img_array[20][2][15] <= img[9087];\
        in_img_array[20][2][16] <= img[9088];\
        in_img_array[20][2][17] <= img[9089];\
        in_img_array[20][3][0] <= img[9090];\
        in_img_array[20][3][1] <= img[9091];\
        in_img_array[20][3][2] <= img[9092];\
        in_img_array[20][3][3] <= img[9093];\
        in_img_array[20][3][4] <= img[9094];\
        in_img_array[20][3][5] <= img[9095];\
        in_img_array[20][3][6] <= img[9096];\
        in_img_array[20][3][7] <= img[9097];\
        in_img_array[20][3][8] <= img[9098];\
        in_img_array[20][3][9] <= img[9099];\
        in_img_array[20][3][10] <= img[9100];\
        in_img_array[20][3][11] <= img[9101];\
        in_img_array[20][3][12] <= img[9102];\
        in_img_array[20][3][13] <= img[9103];\
        in_img_array[20][3][14] <= img[9104];\
        in_img_array[20][3][15] <= img[9105];\
        in_img_array[20][3][16] <= img[9106];\
        in_img_array[20][3][17] <= img[9107];\
        in_img_array[20][4][0] <= img[9108];\
        in_img_array[20][4][1] <= img[9109];\
        in_img_array[20][4][2] <= img[9110];\
        in_img_array[20][4][3] <= img[9111];\
        in_img_array[20][4][4] <= img[9112];\
        in_img_array[20][4][5] <= img[9113];\
        in_img_array[20][4][6] <= img[9114];\
        in_img_array[20][4][7] <= img[9115];\
        in_img_array[20][4][8] <= img[9116];\
        in_img_array[20][4][9] <= img[9117];\
        in_img_array[20][4][10] <= img[9118];\
        in_img_array[20][4][11] <= img[9119];\
        in_img_array[20][4][12] <= img[9120];\
        in_img_array[20][4][13] <= img[9121];\
        in_img_array[20][4][14] <= img[9122];\
        in_img_array[20][4][15] <= img[9123];\
        in_img_array[20][4][16] <= img[9124];\
        in_img_array[20][4][17] <= img[9125];\
        in_img_array[20][5][0] <= img[9126];\
        in_img_array[20][5][1] <= img[9127];\
        in_img_array[20][5][2] <= img[9128];\
        in_img_array[20][5][3] <= img[9129];\
        in_img_array[20][5][4] <= img[9130];\
        in_img_array[20][5][5] <= img[9131];\
        in_img_array[20][5][6] <= img[9132];\
        in_img_array[20][5][7] <= img[9133];\
        in_img_array[20][5][8] <= img[9134];\
        in_img_array[20][5][9] <= img[9135];\
        in_img_array[20][5][10] <= img[9136];\
        in_img_array[20][5][11] <= img[9137];\
        in_img_array[20][5][12] <= img[9138];\
        in_img_array[20][5][13] <= img[9139];\
        in_img_array[20][5][14] <= img[9140];\
        in_img_array[20][5][15] <= img[9141];\
        in_img_array[20][5][16] <= img[9142];\
        in_img_array[20][5][17] <= img[9143];\
        in_img_array[20][6][0] <= img[9144];\
        in_img_array[20][6][1] <= img[9145];\
        in_img_array[20][6][2] <= img[9146];\
        in_img_array[20][6][3] <= img[9147];\
        in_img_array[20][6][4] <= img[9148];\
        in_img_array[20][6][5] <= img[9149];\
        in_img_array[20][6][6] <= img[9150];\
        in_img_array[20][6][7] <= img[9151];\
        in_img_array[20][6][8] <= img[9152];\
        in_img_array[20][6][9] <= img[9153];\
        in_img_array[20][6][10] <= img[9154];\
        in_img_array[20][6][11] <= img[9155];\
        in_img_array[20][6][12] <= img[9156];\
        in_img_array[20][6][13] <= img[9157];\
        in_img_array[20][6][14] <= img[9158];\
        in_img_array[20][6][15] <= img[9159];\
        in_img_array[20][6][16] <= img[9160];\
        in_img_array[20][6][17] <= img[9161];\
        in_img_array[20][7][0] <= img[9162];\
        in_img_array[20][7][1] <= img[9163];\
        in_img_array[20][7][2] <= img[9164];\
        in_img_array[20][7][3] <= img[9165];\
        in_img_array[20][7][4] <= img[9166];\
        in_img_array[20][7][5] <= img[9167];\
        in_img_array[20][7][6] <= img[9168];\
        in_img_array[20][7][7] <= img[9169];\
        in_img_array[20][7][8] <= img[9170];\
        in_img_array[20][7][9] <= img[9171];\
        in_img_array[20][7][10] <= img[9172];\
        in_img_array[20][7][11] <= img[9173];\
        in_img_array[20][7][12] <= img[9174];\
        in_img_array[20][7][13] <= img[9175];\
        in_img_array[20][7][14] <= img[9176];\
        in_img_array[20][7][15] <= img[9177];\
        in_img_array[20][7][16] <= img[9178];\
        in_img_array[20][7][17] <= img[9179];\
        in_img_array[20][8][0] <= img[9180];\
        in_img_array[20][8][1] <= img[9181];\
        in_img_array[20][8][2] <= img[9182];\
        in_img_array[20][8][3] <= img[9183];\
        in_img_array[20][8][4] <= img[9184];\
        in_img_array[20][8][5] <= img[9185];\
        in_img_array[20][8][6] <= img[9186];\
        in_img_array[20][8][7] <= img[9187];\
        in_img_array[20][8][8] <= img[9188];\
        in_img_array[20][8][9] <= img[9189];\
        in_img_array[20][8][10] <= img[9190];\
        in_img_array[20][8][11] <= img[9191];\
        in_img_array[20][8][12] <= img[9192];\
        in_img_array[20][8][13] <= img[9193];\
        in_img_array[20][8][14] <= img[9194];\
        in_img_array[20][8][15] <= img[9195];\
        in_img_array[20][8][16] <= img[9196];\
        in_img_array[20][8][17] <= img[9197];\
        in_img_array[20][9][0] <= img[9198];\
        in_img_array[20][9][1] <= img[9199];\
        in_img_array[20][9][2] <= img[9200];\
        in_img_array[20][9][3] <= img[9201];\
        in_img_array[20][9][4] <= img[9202];\
        in_img_array[20][9][5] <= img[9203];\
        in_img_array[20][9][6] <= img[9204];\
        in_img_array[20][9][7] <= img[9205];\
        in_img_array[20][9][8] <= img[9206];\
        in_img_array[20][9][9] <= img[9207];\
        in_img_array[20][9][10] <= img[9208];\
        in_img_array[20][9][11] <= img[9209];\
        in_img_array[20][9][12] <= img[9210];\
        in_img_array[20][9][13] <= img[9211];\
        in_img_array[20][9][14] <= img[9212];\
        in_img_array[20][9][15] <= img[9213];\
        in_img_array[20][9][16] <= img[9214];\
        in_img_array[20][9][17] <= img[9215];\
        in_img_array[20][10][0] <= img[9216];\
        in_img_array[20][10][1] <= img[9217];\
        in_img_array[20][10][2] <= img[9218];\
        in_img_array[20][10][3] <= img[9219];\
        in_img_array[20][10][4] <= img[9220];\
        in_img_array[20][10][5] <= img[9221];\
        in_img_array[20][10][6] <= img[9222];\
        in_img_array[20][10][7] <= img[9223];\
        in_img_array[20][10][8] <= img[9224];\
        in_img_array[20][10][9] <= img[9225];\
        in_img_array[20][10][10] <= img[9226];\
        in_img_array[20][10][11] <= img[9227];\
        in_img_array[20][10][12] <= img[9228];\
        in_img_array[20][10][13] <= img[9229];\
        in_img_array[20][10][14] <= img[9230];\
        in_img_array[20][10][15] <= img[9231];\
        in_img_array[20][10][16] <= img[9232];\
        in_img_array[20][10][17] <= img[9233];\
        in_img_array[20][11][0] <= img[9234];\
        in_img_array[20][11][1] <= img[9235];\
        in_img_array[20][11][2] <= img[9236];\
        in_img_array[20][11][3] <= img[9237];\
        in_img_array[20][11][4] <= img[9238];\
        in_img_array[20][11][5] <= img[9239];\
        in_img_array[20][11][6] <= img[9240];\
        in_img_array[20][11][7] <= img[9241];\
        in_img_array[20][11][8] <= img[9242];\
        in_img_array[20][11][9] <= img[9243];\
        in_img_array[20][11][10] <= img[9244];\
        in_img_array[20][11][11] <= img[9245];\
        in_img_array[20][11][12] <= img[9246];\
        in_img_array[20][11][13] <= img[9247];\
        in_img_array[20][11][14] <= img[9248];\
        in_img_array[20][11][15] <= img[9249];\
        in_img_array[20][11][16] <= img[9250];\
        in_img_array[20][11][17] <= img[9251];\
        in_img_array[20][12][0] <= img[9252];\
        in_img_array[20][12][1] <= img[9253];\
        in_img_array[20][12][2] <= img[9254];\
        in_img_array[20][12][3] <= img[9255];\
        in_img_array[20][12][4] <= img[9256];\
        in_img_array[20][12][5] <= img[9257];\
        in_img_array[20][12][6] <= img[9258];\
        in_img_array[20][12][7] <= img[9259];\
        in_img_array[20][12][8] <= img[9260];\
        in_img_array[20][12][9] <= img[9261];\
        in_img_array[20][12][10] <= img[9262];\
        in_img_array[20][12][11] <= img[9263];\
        in_img_array[20][12][12] <= img[9264];\
        in_img_array[20][12][13] <= img[9265];\
        in_img_array[20][12][14] <= img[9266];\
        in_img_array[20][12][15] <= img[9267];\
        in_img_array[20][12][16] <= img[9268];\
        in_img_array[20][12][17] <= img[9269];\
        in_img_array[20][13][0] <= img[9270];\
        in_img_array[20][13][1] <= img[9271];\
        in_img_array[20][13][2] <= img[9272];\
        in_img_array[20][13][3] <= img[9273];\
        in_img_array[20][13][4] <= img[9274];\
        in_img_array[20][13][5] <= img[9275];\
        in_img_array[20][13][6] <= img[9276];\
        in_img_array[20][13][7] <= img[9277];\
        in_img_array[20][13][8] <= img[9278];\
        in_img_array[20][13][9] <= img[9279];\
        in_img_array[20][13][10] <= img[9280];\
        in_img_array[20][13][11] <= img[9281];\
        in_img_array[20][13][12] <= img[9282];\
        in_img_array[20][13][13] <= img[9283];\
        in_img_array[20][13][14] <= img[9284];\
        in_img_array[20][13][15] <= img[9285];\
        in_img_array[20][13][16] <= img[9286];\
        in_img_array[20][13][17] <= img[9287];\
        in_img_array[20][14][0] <= img[9288];\
        in_img_array[20][14][1] <= img[9289];\
        in_img_array[20][14][2] <= img[9290];\
        in_img_array[20][14][3] <= img[9291];\
        in_img_array[20][14][4] <= img[9292];\
        in_img_array[20][14][5] <= img[9293];\
        in_img_array[20][14][6] <= img[9294];\
        in_img_array[20][14][7] <= img[9295];\
        in_img_array[20][14][8] <= img[9296];\
        in_img_array[20][14][9] <= img[9297];\
        in_img_array[20][14][10] <= img[9298];\
        in_img_array[20][14][11] <= img[9299];\
        in_img_array[20][14][12] <= img[9300];\
        in_img_array[20][14][13] <= img[9301];\
        in_img_array[20][14][14] <= img[9302];\
        in_img_array[20][14][15] <= img[9303];\
        in_img_array[20][14][16] <= img[9304];\
        in_img_array[20][14][17] <= img[9305];\
        in_img_array[20][15][0] <= img[9306];\
        in_img_array[20][15][1] <= img[9307];\
        in_img_array[20][15][2] <= img[9308];\
        in_img_array[20][15][3] <= img[9309];\
        in_img_array[20][15][4] <= img[9310];\
        in_img_array[20][15][5] <= img[9311];\
        in_img_array[20][15][6] <= img[9312];\
        in_img_array[20][15][7] <= img[9313];\
        in_img_array[20][15][8] <= img[9314];\
        in_img_array[20][15][9] <= img[9315];\
        in_img_array[20][15][10] <= img[9316];\
        in_img_array[20][15][11] <= img[9317];\
        in_img_array[20][15][12] <= img[9318];\
        in_img_array[20][15][13] <= img[9319];\
        in_img_array[20][15][14] <= img[9320];\
        in_img_array[20][15][15] <= img[9321];\
        in_img_array[20][15][16] <= img[9322];\
        in_img_array[20][15][17] <= img[9323];\
        in_img_array[20][16][0] <= img[9324];\
        in_img_array[20][16][1] <= img[9325];\
        in_img_array[20][16][2] <= img[9326];\
        in_img_array[20][16][3] <= img[9327];\
        in_img_array[20][16][4] <= img[9328];\
        in_img_array[20][16][5] <= img[9329];\
        in_img_array[20][16][6] <= img[9330];\
        in_img_array[20][16][7] <= img[9331];\
        in_img_array[20][16][8] <= img[9332];\
        in_img_array[20][16][9] <= img[9333];\
        in_img_array[20][16][10] <= img[9334];\
        in_img_array[20][16][11] <= img[9335];\
        in_img_array[20][16][12] <= img[9336];\
        in_img_array[20][16][13] <= img[9337];\
        in_img_array[20][16][14] <= img[9338];\
        in_img_array[20][16][15] <= img[9339];\
        in_img_array[20][16][16] <= img[9340];\
        in_img_array[20][16][17] <= img[9341];\
        in_img_array[20][17][0] <= img[9342];\
        in_img_array[20][17][1] <= img[9343];\
        in_img_array[20][17][2] <= img[9344];\
        in_img_array[20][17][3] <= img[9345];\
        in_img_array[20][17][4] <= img[9346];\
        in_img_array[20][17][5] <= img[9347];\
        in_img_array[20][17][6] <= img[9348];\
        in_img_array[20][17][7] <= img[9349];\
        in_img_array[20][17][8] <= img[9350];\
        in_img_array[20][17][9] <= img[9351];\
        in_img_array[20][17][10] <= img[9352];\
        in_img_array[20][17][11] <= img[9353];\
        in_img_array[20][17][12] <= img[9354];\
        in_img_array[20][17][13] <= img[9355];\
        in_img_array[20][17][14] <= img[9356];\
        in_img_array[20][17][15] <= img[9357];\
        in_img_array[20][17][16] <= img[9358];\
        in_img_array[20][17][17] <= img[9359];\
        in_img_array[20][18][0] <= img[9360];\
        in_img_array[20][18][1] <= img[9361];\
        in_img_array[20][18][2] <= img[9362];\
        in_img_array[20][18][3] <= img[9363];\
        in_img_array[20][18][4] <= img[9364];\
        in_img_array[20][18][5] <= img[9365];\
        in_img_array[20][18][6] <= img[9366];\
        in_img_array[20][18][7] <= img[9367];\
        in_img_array[20][18][8] <= img[9368];\
        in_img_array[20][18][9] <= img[9369];\
        in_img_array[20][18][10] <= img[9370];\
        in_img_array[20][18][11] <= img[9371];\
        in_img_array[20][18][12] <= img[9372];\
        in_img_array[20][18][13] <= img[9373];\
        in_img_array[20][18][14] <= img[9374];\
        in_img_array[20][18][15] <= img[9375];\
        in_img_array[20][18][16] <= img[9376];\
        in_img_array[20][18][17] <= img[9377];\
        in_img_array[20][19][0] <= img[9378];\
        in_img_array[20][19][1] <= img[9379];\
        in_img_array[20][19][2] <= img[9380];\
        in_img_array[20][19][3] <= img[9381];\
        in_img_array[20][19][4] <= img[9382];\
        in_img_array[20][19][5] <= img[9383];\
        in_img_array[20][19][6] <= img[9384];\
        in_img_array[20][19][7] <= img[9385];\
        in_img_array[20][19][8] <= img[9386];\
        in_img_array[20][19][9] <= img[9387];\
        in_img_array[20][19][10] <= img[9388];\
        in_img_array[20][19][11] <= img[9389];\
        in_img_array[20][19][12] <= img[9390];\
        in_img_array[20][19][13] <= img[9391];\
        in_img_array[20][19][14] <= img[9392];\
        in_img_array[20][19][15] <= img[9393];\
        in_img_array[20][19][16] <= img[9394];\
        in_img_array[20][19][17] <= img[9395];\
        in_img_array[20][20][0] <= img[9396];\
        in_img_array[20][20][1] <= img[9397];\
        in_img_array[20][20][2] <= img[9398];\
        in_img_array[20][20][3] <= img[9399];\
        in_img_array[20][20][4] <= img[9400];\
        in_img_array[20][20][5] <= img[9401];\
        in_img_array[20][20][6] <= img[9402];\
        in_img_array[20][20][7] <= img[9403];\
        in_img_array[20][20][8] <= img[9404];\
        in_img_array[20][20][9] <= img[9405];\
        in_img_array[20][20][10] <= img[9406];\
        in_img_array[20][20][11] <= img[9407];\
        in_img_array[20][20][12] <= img[9408];\
        in_img_array[20][20][13] <= img[9409];\
        in_img_array[20][20][14] <= img[9410];\
        in_img_array[20][20][15] <= img[9411];\
        in_img_array[20][20][16] <= img[9412];\
        in_img_array[20][20][17] <= img[9413];\
        in_img_array[20][21][0] <= img[9414];\
        in_img_array[20][21][1] <= img[9415];\
        in_img_array[20][21][2] <= img[9416];\
        in_img_array[20][21][3] <= img[9417];\
        in_img_array[20][21][4] <= img[9418];\
        in_img_array[20][21][5] <= img[9419];\
        in_img_array[20][21][6] <= img[9420];\
        in_img_array[20][21][7] <= img[9421];\
        in_img_array[20][21][8] <= img[9422];\
        in_img_array[20][21][9] <= img[9423];\
        in_img_array[20][21][10] <= img[9424];\
        in_img_array[20][21][11] <= img[9425];\
        in_img_array[20][21][12] <= img[9426];\
        in_img_array[20][21][13] <= img[9427];\
        in_img_array[20][21][14] <= img[9428];\
        in_img_array[20][21][15] <= img[9429];\
        in_img_array[20][21][16] <= img[9430];\
        in_img_array[20][21][17] <= img[9431];\
        in_img_array[20][22][0] <= img[9432];\
        in_img_array[20][22][1] <= img[9433];\
        in_img_array[20][22][2] <= img[9434];\
        in_img_array[20][22][3] <= img[9435];\
        in_img_array[20][22][4] <= img[9436];\
        in_img_array[20][22][5] <= img[9437];\
        in_img_array[20][22][6] <= img[9438];\
        in_img_array[20][22][7] <= img[9439];\
        in_img_array[20][22][8] <= img[9440];\
        in_img_array[20][22][9] <= img[9441];\
        in_img_array[20][22][10] <= img[9442];\
        in_img_array[20][22][11] <= img[9443];\
        in_img_array[20][22][12] <= img[9444];\
        in_img_array[20][22][13] <= img[9445];\
        in_img_array[20][22][14] <= img[9446];\
        in_img_array[20][22][15] <= img[9447];\
        in_img_array[20][22][16] <= img[9448];\
        in_img_array[20][22][17] <= img[9449];\
        in_img_array[20][23][0] <= img[9450];\
        in_img_array[20][23][1] <= img[9451];\
        in_img_array[20][23][2] <= img[9452];\
        in_img_array[20][23][3] <= img[9453];\
        in_img_array[20][23][4] <= img[9454];\
        in_img_array[20][23][5] <= img[9455];\
        in_img_array[20][23][6] <= img[9456];\
        in_img_array[20][23][7] <= img[9457];\
        in_img_array[20][23][8] <= img[9458];\
        in_img_array[20][23][9] <= img[9459];\
        in_img_array[20][23][10] <= img[9460];\
        in_img_array[20][23][11] <= img[9461];\
        in_img_array[20][23][12] <= img[9462];\
        in_img_array[20][23][13] <= img[9463];\
        in_img_array[20][23][14] <= img[9464];\
        in_img_array[20][23][15] <= img[9465];\
        in_img_array[20][23][16] <= img[9466];\
        in_img_array[20][23][17] <= img[9467];\
        in_img_array[20][24][0] <= img[9468];\
        in_img_array[20][24][1] <= img[9469];\
        in_img_array[20][24][2] <= img[9470];\
        in_img_array[20][24][3] <= img[9471];\
        in_img_array[20][24][4] <= img[9472];\
        in_img_array[20][24][5] <= img[9473];\
        in_img_array[20][24][6] <= img[9474];\
        in_img_array[20][24][7] <= img[9475];\
        in_img_array[20][24][8] <= img[9476];\
        in_img_array[20][24][9] <= img[9477];\
        in_img_array[20][24][10] <= img[9478];\
        in_img_array[20][24][11] <= img[9479];\
        in_img_array[20][24][12] <= img[9480];\
        in_img_array[20][24][13] <= img[9481];\
        in_img_array[20][24][14] <= img[9482];\
        in_img_array[20][24][15] <= img[9483];\
        in_img_array[20][24][16] <= img[9484];\
        in_img_array[20][24][17] <= img[9485];\
        in_img_array[20][25][0] <= img[9486];\
        in_img_array[20][25][1] <= img[9487];\
        in_img_array[20][25][2] <= img[9488];\
        in_img_array[20][25][3] <= img[9489];\
        in_img_array[20][25][4] <= img[9490];\
        in_img_array[20][25][5] <= img[9491];\
        in_img_array[20][25][6] <= img[9492];\
        in_img_array[20][25][7] <= img[9493];\
        in_img_array[20][25][8] <= img[9494];\
        in_img_array[20][25][9] <= img[9495];\
        in_img_array[20][25][10] <= img[9496];\
        in_img_array[20][25][11] <= img[9497];\
        in_img_array[20][25][12] <= img[9498];\
        in_img_array[20][25][13] <= img[9499];\
        in_img_array[20][25][14] <= img[9500];\
        in_img_array[20][25][15] <= img[9501];\
        in_img_array[20][25][16] <= img[9502];\
        in_img_array[20][25][17] <= img[9503];\
        in_img_array[20][26][0] <= img[9504];\
        in_img_array[20][26][1] <= img[9505];\
        in_img_array[20][26][2] <= img[9506];\
        in_img_array[20][26][3] <= img[9507];\
        in_img_array[20][26][4] <= img[9508];\
        in_img_array[20][26][5] <= img[9509];\
        in_img_array[20][26][6] <= img[9510];\
        in_img_array[20][26][7] <= img[9511];\
        in_img_array[20][26][8] <= img[9512];\
        in_img_array[20][26][9] <= img[9513];\
        in_img_array[20][26][10] <= img[9514];\
        in_img_array[20][26][11] <= img[9515];\
        in_img_array[20][26][12] <= img[9516];\
        in_img_array[20][26][13] <= img[9517];\
        in_img_array[20][26][14] <= img[9518];\
        in_img_array[20][26][15] <= img[9519];\
        in_img_array[20][26][16] <= img[9520];\
        in_img_array[20][26][17] <= img[9521];\
        in_img_array[20][27][0] <= img[9522];\
        in_img_array[20][27][1] <= img[9523];\
        in_img_array[20][27][2] <= img[9524];\
        in_img_array[20][27][3] <= img[9525];\
        in_img_array[20][27][4] <= img[9526];\
        in_img_array[20][27][5] <= img[9527];\
        in_img_array[20][27][6] <= img[9528];\
        in_img_array[20][27][7] <= img[9529];\
        in_img_array[20][27][8] <= img[9530];\
        in_img_array[20][27][9] <= img[9531];\
        in_img_array[20][27][10] <= img[9532];\
        in_img_array[20][27][11] <= img[9533];\
        in_img_array[20][27][12] <= img[9534];\
        in_img_array[20][27][13] <= img[9535];\
        in_img_array[20][27][14] <= img[9536];\
        in_img_array[20][27][15] <= img[9537];\
        in_img_array[20][27][16] <= img[9538];\
        in_img_array[20][27][17] <= img[9539];\
        in_img_array[20][28][0] <= img[9540];\
        in_img_array[20][28][1] <= img[9541];\
        in_img_array[20][28][2] <= img[9542];\
        in_img_array[20][28][3] <= img[9543];\
        in_img_array[20][28][4] <= img[9544];\
        in_img_array[20][28][5] <= img[9545];\
        in_img_array[20][28][6] <= img[9546];\
        in_img_array[20][28][7] <= img[9547];\
        in_img_array[20][28][8] <= img[9548];\
        in_img_array[20][28][9] <= img[9549];\
        in_img_array[20][28][10] <= img[9550];\
        in_img_array[20][28][11] <= img[9551];\
        in_img_array[20][28][12] <= img[9552];\
        in_img_array[20][28][13] <= img[9553];\
        in_img_array[20][28][14] <= img[9554];\
        in_img_array[20][28][15] <= img[9555];\
        in_img_array[20][28][16] <= img[9556];\
        in_img_array[20][28][17] <= img[9557];\
        in_img_array[20][29][0] <= img[9558];\
        in_img_array[20][29][1] <= img[9559];\
        in_img_array[20][29][2] <= img[9560];\
        in_img_array[20][29][3] <= img[9561];\
        in_img_array[20][29][4] <= img[9562];\
        in_img_array[20][29][5] <= img[9563];\
        in_img_array[20][29][6] <= img[9564];\
        in_img_array[20][29][7] <= img[9565];\
        in_img_array[20][29][8] <= img[9566];\
        in_img_array[20][29][9] <= img[9567];\
        in_img_array[20][29][10] <= img[9568];\
        in_img_array[20][29][11] <= img[9569];\
        in_img_array[20][29][12] <= img[9570];\
        in_img_array[20][29][13] <= img[9571];\
        in_img_array[20][29][14] <= img[9572];\
        in_img_array[20][29][15] <= img[9573];\
        in_img_array[20][29][16] <= img[9574];\
        in_img_array[20][29][17] <= img[9575];\
        in_img_array[21][2][0] <= img[9576];\
        in_img_array[21][2][1] <= img[9577];\
        in_img_array[21][2][2] <= img[9578];\
        in_img_array[21][2][3] <= img[9579];\
        in_img_array[21][2][4] <= img[9580];\
        in_img_array[21][2][5] <= img[9581];\
        in_img_array[21][2][6] <= img[9582];\
        in_img_array[21][2][7] <= img[9583];\
        in_img_array[21][2][8] <= img[9584];\
        in_img_array[21][2][9] <= img[9585];\
        in_img_array[21][2][10] <= img[9586];\
        in_img_array[21][2][11] <= img[9587];\
        in_img_array[21][2][12] <= img[9588];\
        in_img_array[21][2][13] <= img[9589];\
        in_img_array[21][2][14] <= img[9590];\
        in_img_array[21][2][15] <= img[9591];\
        in_img_array[21][2][16] <= img[9592];\
        in_img_array[21][2][17] <= img[9593];\
        in_img_array[21][3][0] <= img[9594];\
        in_img_array[21][3][1] <= img[9595];\
        in_img_array[21][3][2] <= img[9596];\
        in_img_array[21][3][3] <= img[9597];\
        in_img_array[21][3][4] <= img[9598];\
        in_img_array[21][3][5] <= img[9599];\
        in_img_array[21][3][6] <= img[9600];\
        in_img_array[21][3][7] <= img[9601];\
        in_img_array[21][3][8] <= img[9602];\
        in_img_array[21][3][9] <= img[9603];\
        in_img_array[21][3][10] <= img[9604];\
        in_img_array[21][3][11] <= img[9605];\
        in_img_array[21][3][12] <= img[9606];\
        in_img_array[21][3][13] <= img[9607];\
        in_img_array[21][3][14] <= img[9608];\
        in_img_array[21][3][15] <= img[9609];\
        in_img_array[21][3][16] <= img[9610];\
        in_img_array[21][3][17] <= img[9611];\
        in_img_array[21][4][0] <= img[9612];\
        in_img_array[21][4][1] <= img[9613];\
        in_img_array[21][4][2] <= img[9614];\
        in_img_array[21][4][3] <= img[9615];\
        in_img_array[21][4][4] <= img[9616];\
        in_img_array[21][4][5] <= img[9617];\
        in_img_array[21][4][6] <= img[9618];\
        in_img_array[21][4][7] <= img[9619];\
        in_img_array[21][4][8] <= img[9620];\
        in_img_array[21][4][9] <= img[9621];\
        in_img_array[21][4][10] <= img[9622];\
        in_img_array[21][4][11] <= img[9623];\
        in_img_array[21][4][12] <= img[9624];\
        in_img_array[21][4][13] <= img[9625];\
        in_img_array[21][4][14] <= img[9626];\
        in_img_array[21][4][15] <= img[9627];\
        in_img_array[21][4][16] <= img[9628];\
        in_img_array[21][4][17] <= img[9629];\
        in_img_array[21][5][0] <= img[9630];\
        in_img_array[21][5][1] <= img[9631];\
        in_img_array[21][5][2] <= img[9632];\
        in_img_array[21][5][3] <= img[9633];\
        in_img_array[21][5][4] <= img[9634];\
        in_img_array[21][5][5] <= img[9635];\
        in_img_array[21][5][6] <= img[9636];\
        in_img_array[21][5][7] <= img[9637];\
        in_img_array[21][5][8] <= img[9638];\
        in_img_array[21][5][9] <= img[9639];\
        in_img_array[21][5][10] <= img[9640];\
        in_img_array[21][5][11] <= img[9641];\
        in_img_array[21][5][12] <= img[9642];\
        in_img_array[21][5][13] <= img[9643];\
        in_img_array[21][5][14] <= img[9644];\
        in_img_array[21][5][15] <= img[9645];\
        in_img_array[21][5][16] <= img[9646];\
        in_img_array[21][5][17] <= img[9647];\
        in_img_array[21][6][0] <= img[9648];\
        in_img_array[21][6][1] <= img[9649];\
        in_img_array[21][6][2] <= img[9650];\
        in_img_array[21][6][3] <= img[9651];\
        in_img_array[21][6][4] <= img[9652];\
        in_img_array[21][6][5] <= img[9653];\
        in_img_array[21][6][6] <= img[9654];\
        in_img_array[21][6][7] <= img[9655];\
        in_img_array[21][6][8] <= img[9656];\
        in_img_array[21][6][9] <= img[9657];\
        in_img_array[21][6][10] <= img[9658];\
        in_img_array[21][6][11] <= img[9659];\
        in_img_array[21][6][12] <= img[9660];\
        in_img_array[21][6][13] <= img[9661];\
        in_img_array[21][6][14] <= img[9662];\
        in_img_array[21][6][15] <= img[9663];\
        in_img_array[21][6][16] <= img[9664];\
        in_img_array[21][6][17] <= img[9665];\
        in_img_array[21][7][0] <= img[9666];\
        in_img_array[21][7][1] <= img[9667];\
        in_img_array[21][7][2] <= img[9668];\
        in_img_array[21][7][3] <= img[9669];\
        in_img_array[21][7][4] <= img[9670];\
        in_img_array[21][7][5] <= img[9671];\
        in_img_array[21][7][6] <= img[9672];\
        in_img_array[21][7][7] <= img[9673];\
        in_img_array[21][7][8] <= img[9674];\
        in_img_array[21][7][9] <= img[9675];\
        in_img_array[21][7][10] <= img[9676];\
        in_img_array[21][7][11] <= img[9677];\
        in_img_array[21][7][12] <= img[9678];\
        in_img_array[21][7][13] <= img[9679];\
        in_img_array[21][7][14] <= img[9680];\
        in_img_array[21][7][15] <= img[9681];\
        in_img_array[21][7][16] <= img[9682];\
        in_img_array[21][7][17] <= img[9683];\
        in_img_array[21][8][0] <= img[9684];\
        in_img_array[21][8][1] <= img[9685];\
        in_img_array[21][8][2] <= img[9686];\
        in_img_array[21][8][3] <= img[9687];\
        in_img_array[21][8][4] <= img[9688];\
        in_img_array[21][8][5] <= img[9689];\
        in_img_array[21][8][6] <= img[9690];\
        in_img_array[21][8][7] <= img[9691];\
        in_img_array[21][8][8] <= img[9692];\
        in_img_array[21][8][9] <= img[9693];\
        in_img_array[21][8][10] <= img[9694];\
        in_img_array[21][8][11] <= img[9695];\
        in_img_array[21][8][12] <= img[9696];\
        in_img_array[21][8][13] <= img[9697];\
        in_img_array[21][8][14] <= img[9698];\
        in_img_array[21][8][15] <= img[9699];\
        in_img_array[21][8][16] <= img[9700];\
        in_img_array[21][8][17] <= img[9701];\
        in_img_array[21][9][0] <= img[9702];\
        in_img_array[21][9][1] <= img[9703];\
        in_img_array[21][9][2] <= img[9704];\
        in_img_array[21][9][3] <= img[9705];\
        in_img_array[21][9][4] <= img[9706];\
        in_img_array[21][9][5] <= img[9707];\
        in_img_array[21][9][6] <= img[9708];\
        in_img_array[21][9][7] <= img[9709];\
        in_img_array[21][9][8] <= img[9710];\
        in_img_array[21][9][9] <= img[9711];\
        in_img_array[21][9][10] <= img[9712];\
        in_img_array[21][9][11] <= img[9713];\
        in_img_array[21][9][12] <= img[9714];\
        in_img_array[21][9][13] <= img[9715];\
        in_img_array[21][9][14] <= img[9716];\
        in_img_array[21][9][15] <= img[9717];\
        in_img_array[21][9][16] <= img[9718];\
        in_img_array[21][9][17] <= img[9719];\
        in_img_array[21][10][0] <= img[9720];\
        in_img_array[21][10][1] <= img[9721];\
        in_img_array[21][10][2] <= img[9722];\
        in_img_array[21][10][3] <= img[9723];\
        in_img_array[21][10][4] <= img[9724];\
        in_img_array[21][10][5] <= img[9725];\
        in_img_array[21][10][6] <= img[9726];\
        in_img_array[21][10][7] <= img[9727];\
        in_img_array[21][10][8] <= img[9728];\
        in_img_array[21][10][9] <= img[9729];\
        in_img_array[21][10][10] <= img[9730];\
        in_img_array[21][10][11] <= img[9731];\
        in_img_array[21][10][12] <= img[9732];\
        in_img_array[21][10][13] <= img[9733];\
        in_img_array[21][10][14] <= img[9734];\
        in_img_array[21][10][15] <= img[9735];\
        in_img_array[21][10][16] <= img[9736];\
        in_img_array[21][10][17] <= img[9737];\
        in_img_array[21][11][0] <= img[9738];\
        in_img_array[21][11][1] <= img[9739];\
        in_img_array[21][11][2] <= img[9740];\
        in_img_array[21][11][3] <= img[9741];\
        in_img_array[21][11][4] <= img[9742];\
        in_img_array[21][11][5] <= img[9743];\
        in_img_array[21][11][6] <= img[9744];\
        in_img_array[21][11][7] <= img[9745];\
        in_img_array[21][11][8] <= img[9746];\
        in_img_array[21][11][9] <= img[9747];\
        in_img_array[21][11][10] <= img[9748];\
        in_img_array[21][11][11] <= img[9749];\
        in_img_array[21][11][12] <= img[9750];\
        in_img_array[21][11][13] <= img[9751];\
        in_img_array[21][11][14] <= img[9752];\
        in_img_array[21][11][15] <= img[9753];\
        in_img_array[21][11][16] <= img[9754];\
        in_img_array[21][11][17] <= img[9755];\
        in_img_array[21][12][0] <= img[9756];\
        in_img_array[21][12][1] <= img[9757];\
        in_img_array[21][12][2] <= img[9758];\
        in_img_array[21][12][3] <= img[9759];\
        in_img_array[21][12][4] <= img[9760];\
        in_img_array[21][12][5] <= img[9761];\
        in_img_array[21][12][6] <= img[9762];\
        in_img_array[21][12][7] <= img[9763];\
        in_img_array[21][12][8] <= img[9764];\
        in_img_array[21][12][9] <= img[9765];\
        in_img_array[21][12][10] <= img[9766];\
        in_img_array[21][12][11] <= img[9767];\
        in_img_array[21][12][12] <= img[9768];\
        in_img_array[21][12][13] <= img[9769];\
        in_img_array[21][12][14] <= img[9770];\
        in_img_array[21][12][15] <= img[9771];\
        in_img_array[21][12][16] <= img[9772];\
        in_img_array[21][12][17] <= img[9773];\
        in_img_array[21][13][0] <= img[9774];\
        in_img_array[21][13][1] <= img[9775];\
        in_img_array[21][13][2] <= img[9776];\
        in_img_array[21][13][3] <= img[9777];\
        in_img_array[21][13][4] <= img[9778];\
        in_img_array[21][13][5] <= img[9779];\
        in_img_array[21][13][6] <= img[9780];\
        in_img_array[21][13][7] <= img[9781];\
        in_img_array[21][13][8] <= img[9782];\
        in_img_array[21][13][9] <= img[9783];\
        in_img_array[21][13][10] <= img[9784];\
        in_img_array[21][13][11] <= img[9785];\
        in_img_array[21][13][12] <= img[9786];\
        in_img_array[21][13][13] <= img[9787];\
        in_img_array[21][13][14] <= img[9788];\
        in_img_array[21][13][15] <= img[9789];\
        in_img_array[21][13][16] <= img[9790];\
        in_img_array[21][13][17] <= img[9791];\
        in_img_array[21][14][0] <= img[9792];\
        in_img_array[21][14][1] <= img[9793];\
        in_img_array[21][14][2] <= img[9794];\
        in_img_array[21][14][3] <= img[9795];\
        in_img_array[21][14][4] <= img[9796];\
        in_img_array[21][14][5] <= img[9797];\
        in_img_array[21][14][6] <= img[9798];\
        in_img_array[21][14][7] <= img[9799];\
        in_img_array[21][14][8] <= img[9800];\
        in_img_array[21][14][9] <= img[9801];\
        in_img_array[21][14][10] <= img[9802];\
        in_img_array[21][14][11] <= img[9803];\
        in_img_array[21][14][12] <= img[9804];\
        in_img_array[21][14][13] <= img[9805];\
        in_img_array[21][14][14] <= img[9806];\
        in_img_array[21][14][15] <= img[9807];\
        in_img_array[21][14][16] <= img[9808];\
        in_img_array[21][14][17] <= img[9809];\
        in_img_array[21][15][0] <= img[9810];\
        in_img_array[21][15][1] <= img[9811];\
        in_img_array[21][15][2] <= img[9812];\
        in_img_array[21][15][3] <= img[9813];\
        in_img_array[21][15][4] <= img[9814];\
        in_img_array[21][15][5] <= img[9815];\
        in_img_array[21][15][6] <= img[9816];\
        in_img_array[21][15][7] <= img[9817];\
        in_img_array[21][15][8] <= img[9818];\
        in_img_array[21][15][9] <= img[9819];\
        in_img_array[21][15][10] <= img[9820];\
        in_img_array[21][15][11] <= img[9821];\
        in_img_array[21][15][12] <= img[9822];\
        in_img_array[21][15][13] <= img[9823];\
        in_img_array[21][15][14] <= img[9824];\
        in_img_array[21][15][15] <= img[9825];\
        in_img_array[21][15][16] <= img[9826];\
        in_img_array[21][15][17] <= img[9827];\
        in_img_array[21][16][0] <= img[9828];\
        in_img_array[21][16][1] <= img[9829];\
        in_img_array[21][16][2] <= img[9830];\
        in_img_array[21][16][3] <= img[9831];\
        in_img_array[21][16][4] <= img[9832];\
        in_img_array[21][16][5] <= img[9833];\
        in_img_array[21][16][6] <= img[9834];\
        in_img_array[21][16][7] <= img[9835];\
        in_img_array[21][16][8] <= img[9836];\
        in_img_array[21][16][9] <= img[9837];\
        in_img_array[21][16][10] <= img[9838];\
        in_img_array[21][16][11] <= img[9839];\
        in_img_array[21][16][12] <= img[9840];\
        in_img_array[21][16][13] <= img[9841];\
        in_img_array[21][16][14] <= img[9842];\
        in_img_array[21][16][15] <= img[9843];\
        in_img_array[21][16][16] <= img[9844];\
        in_img_array[21][16][17] <= img[9845];\
        in_img_array[21][17][0] <= img[9846];\
        in_img_array[21][17][1] <= img[9847];\
        in_img_array[21][17][2] <= img[9848];\
        in_img_array[21][17][3] <= img[9849];\
        in_img_array[21][17][4] <= img[9850];\
        in_img_array[21][17][5] <= img[9851];\
        in_img_array[21][17][6] <= img[9852];\
        in_img_array[21][17][7] <= img[9853];\
        in_img_array[21][17][8] <= img[9854];\
        in_img_array[21][17][9] <= img[9855];\
        in_img_array[21][17][10] <= img[9856];\
        in_img_array[21][17][11] <= img[9857];\
        in_img_array[21][17][12] <= img[9858];\
        in_img_array[21][17][13] <= img[9859];\
        in_img_array[21][17][14] <= img[9860];\
        in_img_array[21][17][15] <= img[9861];\
        in_img_array[21][17][16] <= img[9862];\
        in_img_array[21][17][17] <= img[9863];\
        in_img_array[21][18][0] <= img[9864];\
        in_img_array[21][18][1] <= img[9865];\
        in_img_array[21][18][2] <= img[9866];\
        in_img_array[21][18][3] <= img[9867];\
        in_img_array[21][18][4] <= img[9868];\
        in_img_array[21][18][5] <= img[9869];\
        in_img_array[21][18][6] <= img[9870];\
        in_img_array[21][18][7] <= img[9871];\
        in_img_array[21][18][8] <= img[9872];\
        in_img_array[21][18][9] <= img[9873];\
        in_img_array[21][18][10] <= img[9874];\
        in_img_array[21][18][11] <= img[9875];\
        in_img_array[21][18][12] <= img[9876];\
        in_img_array[21][18][13] <= img[9877];\
        in_img_array[21][18][14] <= img[9878];\
        in_img_array[21][18][15] <= img[9879];\
        in_img_array[21][18][16] <= img[9880];\
        in_img_array[21][18][17] <= img[9881];\
        in_img_array[21][19][0] <= img[9882];\
        in_img_array[21][19][1] <= img[9883];\
        in_img_array[21][19][2] <= img[9884];\
        in_img_array[21][19][3] <= img[9885];\
        in_img_array[21][19][4] <= img[9886];\
        in_img_array[21][19][5] <= img[9887];\
        in_img_array[21][19][6] <= img[9888];\
        in_img_array[21][19][7] <= img[9889];\
        in_img_array[21][19][8] <= img[9890];\
        in_img_array[21][19][9] <= img[9891];\
        in_img_array[21][19][10] <= img[9892];\
        in_img_array[21][19][11] <= img[9893];\
        in_img_array[21][19][12] <= img[9894];\
        in_img_array[21][19][13] <= img[9895];\
        in_img_array[21][19][14] <= img[9896];\
        in_img_array[21][19][15] <= img[9897];\
        in_img_array[21][19][16] <= img[9898];\
        in_img_array[21][19][17] <= img[9899];\
        in_img_array[21][20][0] <= img[9900];\
        in_img_array[21][20][1] <= img[9901];\
        in_img_array[21][20][2] <= img[9902];\
        in_img_array[21][20][3] <= img[9903];\
        in_img_array[21][20][4] <= img[9904];\
        in_img_array[21][20][5] <= img[9905];\
        in_img_array[21][20][6] <= img[9906];\
        in_img_array[21][20][7] <= img[9907];\
        in_img_array[21][20][8] <= img[9908];\
        in_img_array[21][20][9] <= img[9909];\
        in_img_array[21][20][10] <= img[9910];\
        in_img_array[21][20][11] <= img[9911];\
        in_img_array[21][20][12] <= img[9912];\
        in_img_array[21][20][13] <= img[9913];\
        in_img_array[21][20][14] <= img[9914];\
        in_img_array[21][20][15] <= img[9915];\
        in_img_array[21][20][16] <= img[9916];\
        in_img_array[21][20][17] <= img[9917];\
        in_img_array[21][21][0] <= img[9918];\
        in_img_array[21][21][1] <= img[9919];\
        in_img_array[21][21][2] <= img[9920];\
        in_img_array[21][21][3] <= img[9921];\
        in_img_array[21][21][4] <= img[9922];\
        in_img_array[21][21][5] <= img[9923];\
        in_img_array[21][21][6] <= img[9924];\
        in_img_array[21][21][7] <= img[9925];\
        in_img_array[21][21][8] <= img[9926];\
        in_img_array[21][21][9] <= img[9927];\
        in_img_array[21][21][10] <= img[9928];\
        in_img_array[21][21][11] <= img[9929];\
        in_img_array[21][21][12] <= img[9930];\
        in_img_array[21][21][13] <= img[9931];\
        in_img_array[21][21][14] <= img[9932];\
        in_img_array[21][21][15] <= img[9933];\
        in_img_array[21][21][16] <= img[9934];\
        in_img_array[21][21][17] <= img[9935];\
        in_img_array[21][22][0] <= img[9936];\
        in_img_array[21][22][1] <= img[9937];\
        in_img_array[21][22][2] <= img[9938];\
        in_img_array[21][22][3] <= img[9939];\
        in_img_array[21][22][4] <= img[9940];\
        in_img_array[21][22][5] <= img[9941];\
        in_img_array[21][22][6] <= img[9942];\
        in_img_array[21][22][7] <= img[9943];\
        in_img_array[21][22][8] <= img[9944];\
        in_img_array[21][22][9] <= img[9945];\
        in_img_array[21][22][10] <= img[9946];\
        in_img_array[21][22][11] <= img[9947];\
        in_img_array[21][22][12] <= img[9948];\
        in_img_array[21][22][13] <= img[9949];\
        in_img_array[21][22][14] <= img[9950];\
        in_img_array[21][22][15] <= img[9951];\
        in_img_array[21][22][16] <= img[9952];\
        in_img_array[21][22][17] <= img[9953];\
        in_img_array[21][23][0] <= img[9954];\
        in_img_array[21][23][1] <= img[9955];\
        in_img_array[21][23][2] <= img[9956];\
        in_img_array[21][23][3] <= img[9957];\
        in_img_array[21][23][4] <= img[9958];\
        in_img_array[21][23][5] <= img[9959];\
        in_img_array[21][23][6] <= img[9960];\
        in_img_array[21][23][7] <= img[9961];\
        in_img_array[21][23][8] <= img[9962];\
        in_img_array[21][23][9] <= img[9963];\
        in_img_array[21][23][10] <= img[9964];\
        in_img_array[21][23][11] <= img[9965];\
        in_img_array[21][23][12] <= img[9966];\
        in_img_array[21][23][13] <= img[9967];\
        in_img_array[21][23][14] <= img[9968];\
        in_img_array[21][23][15] <= img[9969];\
        in_img_array[21][23][16] <= img[9970];\
        in_img_array[21][23][17] <= img[9971];\
        in_img_array[21][24][0] <= img[9972];\
        in_img_array[21][24][1] <= img[9973];\
        in_img_array[21][24][2] <= img[9974];\
        in_img_array[21][24][3] <= img[9975];\
        in_img_array[21][24][4] <= img[9976];\
        in_img_array[21][24][5] <= img[9977];\
        in_img_array[21][24][6] <= img[9978];\
        in_img_array[21][24][7] <= img[9979];\
        in_img_array[21][24][8] <= img[9980];\
        in_img_array[21][24][9] <= img[9981];\
        in_img_array[21][24][10] <= img[9982];\
        in_img_array[21][24][11] <= img[9983];\
        in_img_array[21][24][12] <= img[9984];\
        in_img_array[21][24][13] <= img[9985];\
        in_img_array[21][24][14] <= img[9986];\
        in_img_array[21][24][15] <= img[9987];\
        in_img_array[21][24][16] <= img[9988];\
        in_img_array[21][24][17] <= img[9989];\
        in_img_array[21][25][0] <= img[9990];\
        in_img_array[21][25][1] <= img[9991];\
        in_img_array[21][25][2] <= img[9992];\
        in_img_array[21][25][3] <= img[9993];\
        in_img_array[21][25][4] <= img[9994];\
        in_img_array[21][25][5] <= img[9995];\
        in_img_array[21][25][6] <= img[9996];\
        in_img_array[21][25][7] <= img[9997];\
        in_img_array[21][25][8] <= img[9998];\
        in_img_array[21][25][9] <= img[9999];\
        in_img_array[21][25][10] <= img[10000];\
        in_img_array[21][25][11] <= img[10001];\
        in_img_array[21][25][12] <= img[10002];\
        in_img_array[21][25][13] <= img[10003];\
        in_img_array[21][25][14] <= img[10004];\
        in_img_array[21][25][15] <= img[10005];\
        in_img_array[21][25][16] <= img[10006];\
        in_img_array[21][25][17] <= img[10007];\
        in_img_array[21][26][0] <= img[10008];\
        in_img_array[21][26][1] <= img[10009];\
        in_img_array[21][26][2] <= img[10010];\
        in_img_array[21][26][3] <= img[10011];\
        in_img_array[21][26][4] <= img[10012];\
        in_img_array[21][26][5] <= img[10013];\
        in_img_array[21][26][6] <= img[10014];\
        in_img_array[21][26][7] <= img[10015];\
        in_img_array[21][26][8] <= img[10016];\
        in_img_array[21][26][9] <= img[10017];\
        in_img_array[21][26][10] <= img[10018];\
        in_img_array[21][26][11] <= img[10019];\
        in_img_array[21][26][12] <= img[10020];\
        in_img_array[21][26][13] <= img[10021];\
        in_img_array[21][26][14] <= img[10022];\
        in_img_array[21][26][15] <= img[10023];\
        in_img_array[21][26][16] <= img[10024];\
        in_img_array[21][26][17] <= img[10025];\
        in_img_array[21][27][0] <= img[10026];\
        in_img_array[21][27][1] <= img[10027];\
        in_img_array[21][27][2] <= img[10028];\
        in_img_array[21][27][3] <= img[10029];\
        in_img_array[21][27][4] <= img[10030];\
        in_img_array[21][27][5] <= img[10031];\
        in_img_array[21][27][6] <= img[10032];\
        in_img_array[21][27][7] <= img[10033];\
        in_img_array[21][27][8] <= img[10034];\
        in_img_array[21][27][9] <= img[10035];\
        in_img_array[21][27][10] <= img[10036];\
        in_img_array[21][27][11] <= img[10037];\
        in_img_array[21][27][12] <= img[10038];\
        in_img_array[21][27][13] <= img[10039];\
        in_img_array[21][27][14] <= img[10040];\
        in_img_array[21][27][15] <= img[10041];\
        in_img_array[21][27][16] <= img[10042];\
        in_img_array[21][27][17] <= img[10043];\
        in_img_array[21][28][0] <= img[10044];\
        in_img_array[21][28][1] <= img[10045];\
        in_img_array[21][28][2] <= img[10046];\
        in_img_array[21][28][3] <= img[10047];\
        in_img_array[21][28][4] <= img[10048];\
        in_img_array[21][28][5] <= img[10049];\
        in_img_array[21][28][6] <= img[10050];\
        in_img_array[21][28][7] <= img[10051];\
        in_img_array[21][28][8] <= img[10052];\
        in_img_array[21][28][9] <= img[10053];\
        in_img_array[21][28][10] <= img[10054];\
        in_img_array[21][28][11] <= img[10055];\
        in_img_array[21][28][12] <= img[10056];\
        in_img_array[21][28][13] <= img[10057];\
        in_img_array[21][28][14] <= img[10058];\
        in_img_array[21][28][15] <= img[10059];\
        in_img_array[21][28][16] <= img[10060];\
        in_img_array[21][28][17] <= img[10061];\
        in_img_array[21][29][0] <= img[10062];\
        in_img_array[21][29][1] <= img[10063];\
        in_img_array[21][29][2] <= img[10064];\
        in_img_array[21][29][3] <= img[10065];\
        in_img_array[21][29][4] <= img[10066];\
        in_img_array[21][29][5] <= img[10067];\
        in_img_array[21][29][6] <= img[10068];\
        in_img_array[21][29][7] <= img[10069];\
        in_img_array[21][29][8] <= img[10070];\
        in_img_array[21][29][9] <= img[10071];\
        in_img_array[21][29][10] <= img[10072];\
        in_img_array[21][29][11] <= img[10073];\
        in_img_array[21][29][12] <= img[10074];\
        in_img_array[21][29][13] <= img[10075];\
        in_img_array[21][29][14] <= img[10076];\
        in_img_array[21][29][15] <= img[10077];\
        in_img_array[21][29][16] <= img[10078];\
        in_img_array[21][29][17] <= img[10079];\
        in_img_array[22][2][0] <= img[10080];\
        in_img_array[22][2][1] <= img[10081];\
        in_img_array[22][2][2] <= img[10082];\
        in_img_array[22][2][3] <= img[10083];\
        in_img_array[22][2][4] <= img[10084];\
        in_img_array[22][2][5] <= img[10085];\
        in_img_array[22][2][6] <= img[10086];\
        in_img_array[22][2][7] <= img[10087];\
        in_img_array[22][2][8] <= img[10088];\
        in_img_array[22][2][9] <= img[10089];\
        in_img_array[22][2][10] <= img[10090];\
        in_img_array[22][2][11] <= img[10091];\
        in_img_array[22][2][12] <= img[10092];\
        in_img_array[22][2][13] <= img[10093];\
        in_img_array[22][2][14] <= img[10094];\
        in_img_array[22][2][15] <= img[10095];\
        in_img_array[22][2][16] <= img[10096];\
        in_img_array[22][2][17] <= img[10097];\
        in_img_array[22][3][0] <= img[10098];\
        in_img_array[22][3][1] <= img[10099];\
        in_img_array[22][3][2] <= img[10100];\
        in_img_array[22][3][3] <= img[10101];\
        in_img_array[22][3][4] <= img[10102];\
        in_img_array[22][3][5] <= img[10103];\
        in_img_array[22][3][6] <= img[10104];\
        in_img_array[22][3][7] <= img[10105];\
        in_img_array[22][3][8] <= img[10106];\
        in_img_array[22][3][9] <= img[10107];\
        in_img_array[22][3][10] <= img[10108];\
        in_img_array[22][3][11] <= img[10109];\
        in_img_array[22][3][12] <= img[10110];\
        in_img_array[22][3][13] <= img[10111];\
        in_img_array[22][3][14] <= img[10112];\
        in_img_array[22][3][15] <= img[10113];\
        in_img_array[22][3][16] <= img[10114];\
        in_img_array[22][3][17] <= img[10115];\
        in_img_array[22][4][0] <= img[10116];\
        in_img_array[22][4][1] <= img[10117];\
        in_img_array[22][4][2] <= img[10118];\
        in_img_array[22][4][3] <= img[10119];\
        in_img_array[22][4][4] <= img[10120];\
        in_img_array[22][4][5] <= img[10121];\
        in_img_array[22][4][6] <= img[10122];\
        in_img_array[22][4][7] <= img[10123];\
        in_img_array[22][4][8] <= img[10124];\
        in_img_array[22][4][9] <= img[10125];\
        in_img_array[22][4][10] <= img[10126];\
        in_img_array[22][4][11] <= img[10127];\
        in_img_array[22][4][12] <= img[10128];\
        in_img_array[22][4][13] <= img[10129];\
        in_img_array[22][4][14] <= img[10130];\
        in_img_array[22][4][15] <= img[10131];\
        in_img_array[22][4][16] <= img[10132];\
        in_img_array[22][4][17] <= img[10133];\
        in_img_array[22][5][0] <= img[10134];\
        in_img_array[22][5][1] <= img[10135];\
        in_img_array[22][5][2] <= img[10136];\
        in_img_array[22][5][3] <= img[10137];\
        in_img_array[22][5][4] <= img[10138];\
        in_img_array[22][5][5] <= img[10139];\
        in_img_array[22][5][6] <= img[10140];\
        in_img_array[22][5][7] <= img[10141];\
        in_img_array[22][5][8] <= img[10142];\
        in_img_array[22][5][9] <= img[10143];\
        in_img_array[22][5][10] <= img[10144];\
        in_img_array[22][5][11] <= img[10145];\
        in_img_array[22][5][12] <= img[10146];\
        in_img_array[22][5][13] <= img[10147];\
        in_img_array[22][5][14] <= img[10148];\
        in_img_array[22][5][15] <= img[10149];\
        in_img_array[22][5][16] <= img[10150];\
        in_img_array[22][5][17] <= img[10151];\
        in_img_array[22][6][0] <= img[10152];\
        in_img_array[22][6][1] <= img[10153];\
        in_img_array[22][6][2] <= img[10154];\
        in_img_array[22][6][3] <= img[10155];\
        in_img_array[22][6][4] <= img[10156];\
        in_img_array[22][6][5] <= img[10157];\
        in_img_array[22][6][6] <= img[10158];\
        in_img_array[22][6][7] <= img[10159];\
        in_img_array[22][6][8] <= img[10160];\
        in_img_array[22][6][9] <= img[10161];\
        in_img_array[22][6][10] <= img[10162];\
        in_img_array[22][6][11] <= img[10163];\
        in_img_array[22][6][12] <= img[10164];\
        in_img_array[22][6][13] <= img[10165];\
        in_img_array[22][6][14] <= img[10166];\
        in_img_array[22][6][15] <= img[10167];\
        in_img_array[22][6][16] <= img[10168];\
        in_img_array[22][6][17] <= img[10169];\
        in_img_array[22][7][0] <= img[10170];\
        in_img_array[22][7][1] <= img[10171];\
        in_img_array[22][7][2] <= img[10172];\
        in_img_array[22][7][3] <= img[10173];\
        in_img_array[22][7][4] <= img[10174];\
        in_img_array[22][7][5] <= img[10175];\
        in_img_array[22][7][6] <= img[10176];\
        in_img_array[22][7][7] <= img[10177];\
        in_img_array[22][7][8] <= img[10178];\
        in_img_array[22][7][9] <= img[10179];\
        in_img_array[22][7][10] <= img[10180];\
        in_img_array[22][7][11] <= img[10181];\
        in_img_array[22][7][12] <= img[10182];\
        in_img_array[22][7][13] <= img[10183];\
        in_img_array[22][7][14] <= img[10184];\
        in_img_array[22][7][15] <= img[10185];\
        in_img_array[22][7][16] <= img[10186];\
        in_img_array[22][7][17] <= img[10187];\
        in_img_array[22][8][0] <= img[10188];\
        in_img_array[22][8][1] <= img[10189];\
        in_img_array[22][8][2] <= img[10190];\
        in_img_array[22][8][3] <= img[10191];\
        in_img_array[22][8][4] <= img[10192];\
        in_img_array[22][8][5] <= img[10193];\
        in_img_array[22][8][6] <= img[10194];\
        in_img_array[22][8][7] <= img[10195];\
        in_img_array[22][8][8] <= img[10196];\
        in_img_array[22][8][9] <= img[10197];\
        in_img_array[22][8][10] <= img[10198];\
        in_img_array[22][8][11] <= img[10199];\
        in_img_array[22][8][12] <= img[10200];\
        in_img_array[22][8][13] <= img[10201];\
        in_img_array[22][8][14] <= img[10202];\
        in_img_array[22][8][15] <= img[10203];\
        in_img_array[22][8][16] <= img[10204];\
        in_img_array[22][8][17] <= img[10205];\
        in_img_array[22][9][0] <= img[10206];\
        in_img_array[22][9][1] <= img[10207];\
        in_img_array[22][9][2] <= img[10208];\
        in_img_array[22][9][3] <= img[10209];\
        in_img_array[22][9][4] <= img[10210];\
        in_img_array[22][9][5] <= img[10211];\
        in_img_array[22][9][6] <= img[10212];\
        in_img_array[22][9][7] <= img[10213];\
        in_img_array[22][9][8] <= img[10214];\
        in_img_array[22][9][9] <= img[10215];\
        in_img_array[22][9][10] <= img[10216];\
        in_img_array[22][9][11] <= img[10217];\
        in_img_array[22][9][12] <= img[10218];\
        in_img_array[22][9][13] <= img[10219];\
        in_img_array[22][9][14] <= img[10220];\
        in_img_array[22][9][15] <= img[10221];\
        in_img_array[22][9][16] <= img[10222];\
        in_img_array[22][9][17] <= img[10223];\
        in_img_array[22][10][0] <= img[10224];\
        in_img_array[22][10][1] <= img[10225];\
        in_img_array[22][10][2] <= img[10226];\
        in_img_array[22][10][3] <= img[10227];\
        in_img_array[22][10][4] <= img[10228];\
        in_img_array[22][10][5] <= img[10229];\
        in_img_array[22][10][6] <= img[10230];\
        in_img_array[22][10][7] <= img[10231];\
        in_img_array[22][10][8] <= img[10232];\
        in_img_array[22][10][9] <= img[10233];\
        in_img_array[22][10][10] <= img[10234];\
        in_img_array[22][10][11] <= img[10235];\
        in_img_array[22][10][12] <= img[10236];\
        in_img_array[22][10][13] <= img[10237];\
        in_img_array[22][10][14] <= img[10238];\
        in_img_array[22][10][15] <= img[10239];\
        in_img_array[22][10][16] <= img[10240];\
        in_img_array[22][10][17] <= img[10241];\
        in_img_array[22][11][0] <= img[10242];\
        in_img_array[22][11][1] <= img[10243];\
        in_img_array[22][11][2] <= img[10244];\
        in_img_array[22][11][3] <= img[10245];\
        in_img_array[22][11][4] <= img[10246];\
        in_img_array[22][11][5] <= img[10247];\
        in_img_array[22][11][6] <= img[10248];\
        in_img_array[22][11][7] <= img[10249];\
        in_img_array[22][11][8] <= img[10250];\
        in_img_array[22][11][9] <= img[10251];\
        in_img_array[22][11][10] <= img[10252];\
        in_img_array[22][11][11] <= img[10253];\
        in_img_array[22][11][12] <= img[10254];\
        in_img_array[22][11][13] <= img[10255];\
        in_img_array[22][11][14] <= img[10256];\
        in_img_array[22][11][15] <= img[10257];\
        in_img_array[22][11][16] <= img[10258];\
        in_img_array[22][11][17] <= img[10259];\
        in_img_array[22][12][0] <= img[10260];\
        in_img_array[22][12][1] <= img[10261];\
        in_img_array[22][12][2] <= img[10262];\
        in_img_array[22][12][3] <= img[10263];\
        in_img_array[22][12][4] <= img[10264];\
        in_img_array[22][12][5] <= img[10265];\
        in_img_array[22][12][6] <= img[10266];\
        in_img_array[22][12][7] <= img[10267];\
        in_img_array[22][12][8] <= img[10268];\
        in_img_array[22][12][9] <= img[10269];\
        in_img_array[22][12][10] <= img[10270];\
        in_img_array[22][12][11] <= img[10271];\
        in_img_array[22][12][12] <= img[10272];\
        in_img_array[22][12][13] <= img[10273];\
        in_img_array[22][12][14] <= img[10274];\
        in_img_array[22][12][15] <= img[10275];\
        in_img_array[22][12][16] <= img[10276];\
        in_img_array[22][12][17] <= img[10277];\
        in_img_array[22][13][0] <= img[10278];\
        in_img_array[22][13][1] <= img[10279];\
        in_img_array[22][13][2] <= img[10280];\
        in_img_array[22][13][3] <= img[10281];\
        in_img_array[22][13][4] <= img[10282];\
        in_img_array[22][13][5] <= img[10283];\
        in_img_array[22][13][6] <= img[10284];\
        in_img_array[22][13][7] <= img[10285];\
        in_img_array[22][13][8] <= img[10286];\
        in_img_array[22][13][9] <= img[10287];\
        in_img_array[22][13][10] <= img[10288];\
        in_img_array[22][13][11] <= img[10289];\
        in_img_array[22][13][12] <= img[10290];\
        in_img_array[22][13][13] <= img[10291];\
        in_img_array[22][13][14] <= img[10292];\
        in_img_array[22][13][15] <= img[10293];\
        in_img_array[22][13][16] <= img[10294];\
        in_img_array[22][13][17] <= img[10295];\
        in_img_array[22][14][0] <= img[10296];\
        in_img_array[22][14][1] <= img[10297];\
        in_img_array[22][14][2] <= img[10298];\
        in_img_array[22][14][3] <= img[10299];\
        in_img_array[22][14][4] <= img[10300];\
        in_img_array[22][14][5] <= img[10301];\
        in_img_array[22][14][6] <= img[10302];\
        in_img_array[22][14][7] <= img[10303];\
        in_img_array[22][14][8] <= img[10304];\
        in_img_array[22][14][9] <= img[10305];\
        in_img_array[22][14][10] <= img[10306];\
        in_img_array[22][14][11] <= img[10307];\
        in_img_array[22][14][12] <= img[10308];\
        in_img_array[22][14][13] <= img[10309];\
        in_img_array[22][14][14] <= img[10310];\
        in_img_array[22][14][15] <= img[10311];\
        in_img_array[22][14][16] <= img[10312];\
        in_img_array[22][14][17] <= img[10313];\
        in_img_array[22][15][0] <= img[10314];\
        in_img_array[22][15][1] <= img[10315];\
        in_img_array[22][15][2] <= img[10316];\
        in_img_array[22][15][3] <= img[10317];\
        in_img_array[22][15][4] <= img[10318];\
        in_img_array[22][15][5] <= img[10319];\
        in_img_array[22][15][6] <= img[10320];\
        in_img_array[22][15][7] <= img[10321];\
        in_img_array[22][15][8] <= img[10322];\
        in_img_array[22][15][9] <= img[10323];\
        in_img_array[22][15][10] <= img[10324];\
        in_img_array[22][15][11] <= img[10325];\
        in_img_array[22][15][12] <= img[10326];\
        in_img_array[22][15][13] <= img[10327];\
        in_img_array[22][15][14] <= img[10328];\
        in_img_array[22][15][15] <= img[10329];\
        in_img_array[22][15][16] <= img[10330];\
        in_img_array[22][15][17] <= img[10331];\
        in_img_array[22][16][0] <= img[10332];\
        in_img_array[22][16][1] <= img[10333];\
        in_img_array[22][16][2] <= img[10334];\
        in_img_array[22][16][3] <= img[10335];\
        in_img_array[22][16][4] <= img[10336];\
        in_img_array[22][16][5] <= img[10337];\
        in_img_array[22][16][6] <= img[10338];\
        in_img_array[22][16][7] <= img[10339];\
        in_img_array[22][16][8] <= img[10340];\
        in_img_array[22][16][9] <= img[10341];\
        in_img_array[22][16][10] <= img[10342];\
        in_img_array[22][16][11] <= img[10343];\
        in_img_array[22][16][12] <= img[10344];\
        in_img_array[22][16][13] <= img[10345];\
        in_img_array[22][16][14] <= img[10346];\
        in_img_array[22][16][15] <= img[10347];\
        in_img_array[22][16][16] <= img[10348];\
        in_img_array[22][16][17] <= img[10349];\
        in_img_array[22][17][0] <= img[10350];\
        in_img_array[22][17][1] <= img[10351];\
        in_img_array[22][17][2] <= img[10352];\
        in_img_array[22][17][3] <= img[10353];\
        in_img_array[22][17][4] <= img[10354];\
        in_img_array[22][17][5] <= img[10355];\
        in_img_array[22][17][6] <= img[10356];\
        in_img_array[22][17][7] <= img[10357];\
        in_img_array[22][17][8] <= img[10358];\
        in_img_array[22][17][9] <= img[10359];\
        in_img_array[22][17][10] <= img[10360];\
        in_img_array[22][17][11] <= img[10361];\
        in_img_array[22][17][12] <= img[10362];\
        in_img_array[22][17][13] <= img[10363];\
        in_img_array[22][17][14] <= img[10364];\
        in_img_array[22][17][15] <= img[10365];\
        in_img_array[22][17][16] <= img[10366];\
        in_img_array[22][17][17] <= img[10367];\
        in_img_array[22][18][0] <= img[10368];\
        in_img_array[22][18][1] <= img[10369];\
        in_img_array[22][18][2] <= img[10370];\
        in_img_array[22][18][3] <= img[10371];\
        in_img_array[22][18][4] <= img[10372];\
        in_img_array[22][18][5] <= img[10373];\
        in_img_array[22][18][6] <= img[10374];\
        in_img_array[22][18][7] <= img[10375];\
        in_img_array[22][18][8] <= img[10376];\
        in_img_array[22][18][9] <= img[10377];\
        in_img_array[22][18][10] <= img[10378];\
        in_img_array[22][18][11] <= img[10379];\
        in_img_array[22][18][12] <= img[10380];\
        in_img_array[22][18][13] <= img[10381];\
        in_img_array[22][18][14] <= img[10382];\
        in_img_array[22][18][15] <= img[10383];\
        in_img_array[22][18][16] <= img[10384];\
        in_img_array[22][18][17] <= img[10385];\
        in_img_array[22][19][0] <= img[10386];\
        in_img_array[22][19][1] <= img[10387];\
        in_img_array[22][19][2] <= img[10388];\
        in_img_array[22][19][3] <= img[10389];\
        in_img_array[22][19][4] <= img[10390];\
        in_img_array[22][19][5] <= img[10391];\
        in_img_array[22][19][6] <= img[10392];\
        in_img_array[22][19][7] <= img[10393];\
        in_img_array[22][19][8] <= img[10394];\
        in_img_array[22][19][9] <= img[10395];\
        in_img_array[22][19][10] <= img[10396];\
        in_img_array[22][19][11] <= img[10397];\
        in_img_array[22][19][12] <= img[10398];\
        in_img_array[22][19][13] <= img[10399];\
        in_img_array[22][19][14] <= img[10400];\
        in_img_array[22][19][15] <= img[10401];\
        in_img_array[22][19][16] <= img[10402];\
        in_img_array[22][19][17] <= img[10403];\
        in_img_array[22][20][0] <= img[10404];\
        in_img_array[22][20][1] <= img[10405];\
        in_img_array[22][20][2] <= img[10406];\
        in_img_array[22][20][3] <= img[10407];\
        in_img_array[22][20][4] <= img[10408];\
        in_img_array[22][20][5] <= img[10409];\
        in_img_array[22][20][6] <= img[10410];\
        in_img_array[22][20][7] <= img[10411];\
        in_img_array[22][20][8] <= img[10412];\
        in_img_array[22][20][9] <= img[10413];\
        in_img_array[22][20][10] <= img[10414];\
        in_img_array[22][20][11] <= img[10415];\
        in_img_array[22][20][12] <= img[10416];\
        in_img_array[22][20][13] <= img[10417];\
        in_img_array[22][20][14] <= img[10418];\
        in_img_array[22][20][15] <= img[10419];\
        in_img_array[22][20][16] <= img[10420];\
        in_img_array[22][20][17] <= img[10421];\
        in_img_array[22][21][0] <= img[10422];\
        in_img_array[22][21][1] <= img[10423];\
        in_img_array[22][21][2] <= img[10424];\
        in_img_array[22][21][3] <= img[10425];\
        in_img_array[22][21][4] <= img[10426];\
        in_img_array[22][21][5] <= img[10427];\
        in_img_array[22][21][6] <= img[10428];\
        in_img_array[22][21][7] <= img[10429];\
        in_img_array[22][21][8] <= img[10430];\
        in_img_array[22][21][9] <= img[10431];\
        in_img_array[22][21][10] <= img[10432];\
        in_img_array[22][21][11] <= img[10433];\
        in_img_array[22][21][12] <= img[10434];\
        in_img_array[22][21][13] <= img[10435];\
        in_img_array[22][21][14] <= img[10436];\
        in_img_array[22][21][15] <= img[10437];\
        in_img_array[22][21][16] <= img[10438];\
        in_img_array[22][21][17] <= img[10439];\
        in_img_array[22][22][0] <= img[10440];\
        in_img_array[22][22][1] <= img[10441];\
        in_img_array[22][22][2] <= img[10442];\
        in_img_array[22][22][3] <= img[10443];\
        in_img_array[22][22][4] <= img[10444];\
        in_img_array[22][22][5] <= img[10445];\
        in_img_array[22][22][6] <= img[10446];\
        in_img_array[22][22][7] <= img[10447];\
        in_img_array[22][22][8] <= img[10448];\
        in_img_array[22][22][9] <= img[10449];\
        in_img_array[22][22][10] <= img[10450];\
        in_img_array[22][22][11] <= img[10451];\
        in_img_array[22][22][12] <= img[10452];\
        in_img_array[22][22][13] <= img[10453];\
        in_img_array[22][22][14] <= img[10454];\
        in_img_array[22][22][15] <= img[10455];\
        in_img_array[22][22][16] <= img[10456];\
        in_img_array[22][22][17] <= img[10457];\
        in_img_array[22][23][0] <= img[10458];\
        in_img_array[22][23][1] <= img[10459];\
        in_img_array[22][23][2] <= img[10460];\
        in_img_array[22][23][3] <= img[10461];\
        in_img_array[22][23][4] <= img[10462];\
        in_img_array[22][23][5] <= img[10463];\
        in_img_array[22][23][6] <= img[10464];\
        in_img_array[22][23][7] <= img[10465];\
        in_img_array[22][23][8] <= img[10466];\
        in_img_array[22][23][9] <= img[10467];\
        in_img_array[22][23][10] <= img[10468];\
        in_img_array[22][23][11] <= img[10469];\
        in_img_array[22][23][12] <= img[10470];\
        in_img_array[22][23][13] <= img[10471];\
        in_img_array[22][23][14] <= img[10472];\
        in_img_array[22][23][15] <= img[10473];\
        in_img_array[22][23][16] <= img[10474];\
        in_img_array[22][23][17] <= img[10475];\
        in_img_array[22][24][0] <= img[10476];\
        in_img_array[22][24][1] <= img[10477];\
        in_img_array[22][24][2] <= img[10478];\
        in_img_array[22][24][3] <= img[10479];\
        in_img_array[22][24][4] <= img[10480];\
        in_img_array[22][24][5] <= img[10481];\
        in_img_array[22][24][6] <= img[10482];\
        in_img_array[22][24][7] <= img[10483];\
        in_img_array[22][24][8] <= img[10484];\
        in_img_array[22][24][9] <= img[10485];\
        in_img_array[22][24][10] <= img[10486];\
        in_img_array[22][24][11] <= img[10487];\
        in_img_array[22][24][12] <= img[10488];\
        in_img_array[22][24][13] <= img[10489];\
        in_img_array[22][24][14] <= img[10490];\
        in_img_array[22][24][15] <= img[10491];\
        in_img_array[22][24][16] <= img[10492];\
        in_img_array[22][24][17] <= img[10493];\
        in_img_array[22][25][0] <= img[10494];\
        in_img_array[22][25][1] <= img[10495];\
        in_img_array[22][25][2] <= img[10496];\
        in_img_array[22][25][3] <= img[10497];\
        in_img_array[22][25][4] <= img[10498];\
        in_img_array[22][25][5] <= img[10499];\
        in_img_array[22][25][6] <= img[10500];\
        in_img_array[22][25][7] <= img[10501];\
        in_img_array[22][25][8] <= img[10502];\
        in_img_array[22][25][9] <= img[10503];\
        in_img_array[22][25][10] <= img[10504];\
        in_img_array[22][25][11] <= img[10505];\
        in_img_array[22][25][12] <= img[10506];\
        in_img_array[22][25][13] <= img[10507];\
        in_img_array[22][25][14] <= img[10508];\
        in_img_array[22][25][15] <= img[10509];\
        in_img_array[22][25][16] <= img[10510];\
        in_img_array[22][25][17] <= img[10511];\
        in_img_array[22][26][0] <= img[10512];\
        in_img_array[22][26][1] <= img[10513];\
        in_img_array[22][26][2] <= img[10514];\
        in_img_array[22][26][3] <= img[10515];\
        in_img_array[22][26][4] <= img[10516];\
        in_img_array[22][26][5] <= img[10517];\
        in_img_array[22][26][6] <= img[10518];\
        in_img_array[22][26][7] <= img[10519];\
        in_img_array[22][26][8] <= img[10520];\
        in_img_array[22][26][9] <= img[10521];\
        in_img_array[22][26][10] <= img[10522];\
        in_img_array[22][26][11] <= img[10523];\
        in_img_array[22][26][12] <= img[10524];\
        in_img_array[22][26][13] <= img[10525];\
        in_img_array[22][26][14] <= img[10526];\
        in_img_array[22][26][15] <= img[10527];\
        in_img_array[22][26][16] <= img[10528];\
        in_img_array[22][26][17] <= img[10529];\
        in_img_array[22][27][0] <= img[10530];\
        in_img_array[22][27][1] <= img[10531];\
        in_img_array[22][27][2] <= img[10532];\
        in_img_array[22][27][3] <= img[10533];\
        in_img_array[22][27][4] <= img[10534];\
        in_img_array[22][27][5] <= img[10535];\
        in_img_array[22][27][6] <= img[10536];\
        in_img_array[22][27][7] <= img[10537];\
        in_img_array[22][27][8] <= img[10538];\
        in_img_array[22][27][9] <= img[10539];\
        in_img_array[22][27][10] <= img[10540];\
        in_img_array[22][27][11] <= img[10541];\
        in_img_array[22][27][12] <= img[10542];\
        in_img_array[22][27][13] <= img[10543];\
        in_img_array[22][27][14] <= img[10544];\
        in_img_array[22][27][15] <= img[10545];\
        in_img_array[22][27][16] <= img[10546];\
        in_img_array[22][27][17] <= img[10547];\
        in_img_array[22][28][0] <= img[10548];\
        in_img_array[22][28][1] <= img[10549];\
        in_img_array[22][28][2] <= img[10550];\
        in_img_array[22][28][3] <= img[10551];\
        in_img_array[22][28][4] <= img[10552];\
        in_img_array[22][28][5] <= img[10553];\
        in_img_array[22][28][6] <= img[10554];\
        in_img_array[22][28][7] <= img[10555];\
        in_img_array[22][28][8] <= img[10556];\
        in_img_array[22][28][9] <= img[10557];\
        in_img_array[22][28][10] <= img[10558];\
        in_img_array[22][28][11] <= img[10559];\
        in_img_array[22][28][12] <= img[10560];\
        in_img_array[22][28][13] <= img[10561];\
        in_img_array[22][28][14] <= img[10562];\
        in_img_array[22][28][15] <= img[10563];\
        in_img_array[22][28][16] <= img[10564];\
        in_img_array[22][28][17] <= img[10565];\
        in_img_array[22][29][0] <= img[10566];\
        in_img_array[22][29][1] <= img[10567];\
        in_img_array[22][29][2] <= img[10568];\
        in_img_array[22][29][3] <= img[10569];\
        in_img_array[22][29][4] <= img[10570];\
        in_img_array[22][29][5] <= img[10571];\
        in_img_array[22][29][6] <= img[10572];\
        in_img_array[22][29][7] <= img[10573];\
        in_img_array[22][29][8] <= img[10574];\
        in_img_array[22][29][9] <= img[10575];\
        in_img_array[22][29][10] <= img[10576];\
        in_img_array[22][29][11] <= img[10577];\
        in_img_array[22][29][12] <= img[10578];\
        in_img_array[22][29][13] <= img[10579];\
        in_img_array[22][29][14] <= img[10580];\
        in_img_array[22][29][15] <= img[10581];\
        in_img_array[22][29][16] <= img[10582];\
        in_img_array[22][29][17] <= img[10583];\
        in_img_array[23][2][0] <= img[10584];\
        in_img_array[23][2][1] <= img[10585];\
        in_img_array[23][2][2] <= img[10586];\
        in_img_array[23][2][3] <= img[10587];\
        in_img_array[23][2][4] <= img[10588];\
        in_img_array[23][2][5] <= img[10589];\
        in_img_array[23][2][6] <= img[10590];\
        in_img_array[23][2][7] <= img[10591];\
        in_img_array[23][2][8] <= img[10592];\
        in_img_array[23][2][9] <= img[10593];\
        in_img_array[23][2][10] <= img[10594];\
        in_img_array[23][2][11] <= img[10595];\
        in_img_array[23][2][12] <= img[10596];\
        in_img_array[23][2][13] <= img[10597];\
        in_img_array[23][2][14] <= img[10598];\
        in_img_array[23][2][15] <= img[10599];\
        in_img_array[23][2][16] <= img[10600];\
        in_img_array[23][2][17] <= img[10601];\
        in_img_array[23][3][0] <= img[10602];\
        in_img_array[23][3][1] <= img[10603];\
        in_img_array[23][3][2] <= img[10604];\
        in_img_array[23][3][3] <= img[10605];\
        in_img_array[23][3][4] <= img[10606];\
        in_img_array[23][3][5] <= img[10607];\
        in_img_array[23][3][6] <= img[10608];\
        in_img_array[23][3][7] <= img[10609];\
        in_img_array[23][3][8] <= img[10610];\
        in_img_array[23][3][9] <= img[10611];\
        in_img_array[23][3][10] <= img[10612];\
        in_img_array[23][3][11] <= img[10613];\
        in_img_array[23][3][12] <= img[10614];\
        in_img_array[23][3][13] <= img[10615];\
        in_img_array[23][3][14] <= img[10616];\
        in_img_array[23][3][15] <= img[10617];\
        in_img_array[23][3][16] <= img[10618];\
        in_img_array[23][3][17] <= img[10619];\
        in_img_array[23][4][0] <= img[10620];\
        in_img_array[23][4][1] <= img[10621];\
        in_img_array[23][4][2] <= img[10622];\
        in_img_array[23][4][3] <= img[10623];\
        in_img_array[23][4][4] <= img[10624];\
        in_img_array[23][4][5] <= img[10625];\
        in_img_array[23][4][6] <= img[10626];\
        in_img_array[23][4][7] <= img[10627];\
        in_img_array[23][4][8] <= img[10628];\
        in_img_array[23][4][9] <= img[10629];\
        in_img_array[23][4][10] <= img[10630];\
        in_img_array[23][4][11] <= img[10631];\
        in_img_array[23][4][12] <= img[10632];\
        in_img_array[23][4][13] <= img[10633];\
        in_img_array[23][4][14] <= img[10634];\
        in_img_array[23][4][15] <= img[10635];\
        in_img_array[23][4][16] <= img[10636];\
        in_img_array[23][4][17] <= img[10637];\
        in_img_array[23][5][0] <= img[10638];\
        in_img_array[23][5][1] <= img[10639];\
        in_img_array[23][5][2] <= img[10640];\
        in_img_array[23][5][3] <= img[10641];\
        in_img_array[23][5][4] <= img[10642];\
        in_img_array[23][5][5] <= img[10643];\
        in_img_array[23][5][6] <= img[10644];\
        in_img_array[23][5][7] <= img[10645];\
        in_img_array[23][5][8] <= img[10646];\
        in_img_array[23][5][9] <= img[10647];\
        in_img_array[23][5][10] <= img[10648];\
        in_img_array[23][5][11] <= img[10649];\
        in_img_array[23][5][12] <= img[10650];\
        in_img_array[23][5][13] <= img[10651];\
        in_img_array[23][5][14] <= img[10652];\
        in_img_array[23][5][15] <= img[10653];\
        in_img_array[23][5][16] <= img[10654];\
        in_img_array[23][5][17] <= img[10655];\
        in_img_array[23][6][0] <= img[10656];\
        in_img_array[23][6][1] <= img[10657];\
        in_img_array[23][6][2] <= img[10658];\
        in_img_array[23][6][3] <= img[10659];\
        in_img_array[23][6][4] <= img[10660];\
        in_img_array[23][6][5] <= img[10661];\
        in_img_array[23][6][6] <= img[10662];\
        in_img_array[23][6][7] <= img[10663];\
        in_img_array[23][6][8] <= img[10664];\
        in_img_array[23][6][9] <= img[10665];\
        in_img_array[23][6][10] <= img[10666];\
        in_img_array[23][6][11] <= img[10667];\
        in_img_array[23][6][12] <= img[10668];\
        in_img_array[23][6][13] <= img[10669];\
        in_img_array[23][6][14] <= img[10670];\
        in_img_array[23][6][15] <= img[10671];\
        in_img_array[23][6][16] <= img[10672];\
        in_img_array[23][6][17] <= img[10673];\
        in_img_array[23][7][0] <= img[10674];\
        in_img_array[23][7][1] <= img[10675];\
        in_img_array[23][7][2] <= img[10676];\
        in_img_array[23][7][3] <= img[10677];\
        in_img_array[23][7][4] <= img[10678];\
        in_img_array[23][7][5] <= img[10679];\
        in_img_array[23][7][6] <= img[10680];\
        in_img_array[23][7][7] <= img[10681];\
        in_img_array[23][7][8] <= img[10682];\
        in_img_array[23][7][9] <= img[10683];\
        in_img_array[23][7][10] <= img[10684];\
        in_img_array[23][7][11] <= img[10685];\
        in_img_array[23][7][12] <= img[10686];\
        in_img_array[23][7][13] <= img[10687];\
        in_img_array[23][7][14] <= img[10688];\
        in_img_array[23][7][15] <= img[10689];\
        in_img_array[23][7][16] <= img[10690];\
        in_img_array[23][7][17] <= img[10691];\
        in_img_array[23][8][0] <= img[10692];\
        in_img_array[23][8][1] <= img[10693];\
        in_img_array[23][8][2] <= img[10694];\
        in_img_array[23][8][3] <= img[10695];\
        in_img_array[23][8][4] <= img[10696];\
        in_img_array[23][8][5] <= img[10697];\
        in_img_array[23][8][6] <= img[10698];\
        in_img_array[23][8][7] <= img[10699];\
        in_img_array[23][8][8] <= img[10700];\
        in_img_array[23][8][9] <= img[10701];\
        in_img_array[23][8][10] <= img[10702];\
        in_img_array[23][8][11] <= img[10703];\
        in_img_array[23][8][12] <= img[10704];\
        in_img_array[23][8][13] <= img[10705];\
        in_img_array[23][8][14] <= img[10706];\
        in_img_array[23][8][15] <= img[10707];\
        in_img_array[23][8][16] <= img[10708];\
        in_img_array[23][8][17] <= img[10709];\
        in_img_array[23][9][0] <= img[10710];\
        in_img_array[23][9][1] <= img[10711];\
        in_img_array[23][9][2] <= img[10712];\
        in_img_array[23][9][3] <= img[10713];\
        in_img_array[23][9][4] <= img[10714];\
        in_img_array[23][9][5] <= img[10715];\
        in_img_array[23][9][6] <= img[10716];\
        in_img_array[23][9][7] <= img[10717];\
        in_img_array[23][9][8] <= img[10718];\
        in_img_array[23][9][9] <= img[10719];\
        in_img_array[23][9][10] <= img[10720];\
        in_img_array[23][9][11] <= img[10721];\
        in_img_array[23][9][12] <= img[10722];\
        in_img_array[23][9][13] <= img[10723];\
        in_img_array[23][9][14] <= img[10724];\
        in_img_array[23][9][15] <= img[10725];\
        in_img_array[23][9][16] <= img[10726];\
        in_img_array[23][9][17] <= img[10727];\
        in_img_array[23][10][0] <= img[10728];\
        in_img_array[23][10][1] <= img[10729];\
        in_img_array[23][10][2] <= img[10730];\
        in_img_array[23][10][3] <= img[10731];\
        in_img_array[23][10][4] <= img[10732];\
        in_img_array[23][10][5] <= img[10733];\
        in_img_array[23][10][6] <= img[10734];\
        in_img_array[23][10][7] <= img[10735];\
        in_img_array[23][10][8] <= img[10736];\
        in_img_array[23][10][9] <= img[10737];\
        in_img_array[23][10][10] <= img[10738];\
        in_img_array[23][10][11] <= img[10739];\
        in_img_array[23][10][12] <= img[10740];\
        in_img_array[23][10][13] <= img[10741];\
        in_img_array[23][10][14] <= img[10742];\
        in_img_array[23][10][15] <= img[10743];\
        in_img_array[23][10][16] <= img[10744];\
        in_img_array[23][10][17] <= img[10745];\
        in_img_array[23][11][0] <= img[10746];\
        in_img_array[23][11][1] <= img[10747];\
        in_img_array[23][11][2] <= img[10748];\
        in_img_array[23][11][3] <= img[10749];\
        in_img_array[23][11][4] <= img[10750];\
        in_img_array[23][11][5] <= img[10751];\
        in_img_array[23][11][6] <= img[10752];\
        in_img_array[23][11][7] <= img[10753];\
        in_img_array[23][11][8] <= img[10754];\
        in_img_array[23][11][9] <= img[10755];\
        in_img_array[23][11][10] <= img[10756];\
        in_img_array[23][11][11] <= img[10757];\
        in_img_array[23][11][12] <= img[10758];\
        in_img_array[23][11][13] <= img[10759];\
        in_img_array[23][11][14] <= img[10760];\
        in_img_array[23][11][15] <= img[10761];\
        in_img_array[23][11][16] <= img[10762];\
        in_img_array[23][11][17] <= img[10763];\
        in_img_array[23][12][0] <= img[10764];\
        in_img_array[23][12][1] <= img[10765];\
        in_img_array[23][12][2] <= img[10766];\
        in_img_array[23][12][3] <= img[10767];\
        in_img_array[23][12][4] <= img[10768];\
        in_img_array[23][12][5] <= img[10769];\
        in_img_array[23][12][6] <= img[10770];\
        in_img_array[23][12][7] <= img[10771];\
        in_img_array[23][12][8] <= img[10772];\
        in_img_array[23][12][9] <= img[10773];\
        in_img_array[23][12][10] <= img[10774];\
        in_img_array[23][12][11] <= img[10775];\
        in_img_array[23][12][12] <= img[10776];\
        in_img_array[23][12][13] <= img[10777];\
        in_img_array[23][12][14] <= img[10778];\
        in_img_array[23][12][15] <= img[10779];\
        in_img_array[23][12][16] <= img[10780];\
        in_img_array[23][12][17] <= img[10781];\
        in_img_array[23][13][0] <= img[10782];\
        in_img_array[23][13][1] <= img[10783];\
        in_img_array[23][13][2] <= img[10784];\
        in_img_array[23][13][3] <= img[10785];\
        in_img_array[23][13][4] <= img[10786];\
        in_img_array[23][13][5] <= img[10787];\
        in_img_array[23][13][6] <= img[10788];\
        in_img_array[23][13][7] <= img[10789];\
        in_img_array[23][13][8] <= img[10790];\
        in_img_array[23][13][9] <= img[10791];\
        in_img_array[23][13][10] <= img[10792];\
        in_img_array[23][13][11] <= img[10793];\
        in_img_array[23][13][12] <= img[10794];\
        in_img_array[23][13][13] <= img[10795];\
        in_img_array[23][13][14] <= img[10796];\
        in_img_array[23][13][15] <= img[10797];\
        in_img_array[23][13][16] <= img[10798];\
        in_img_array[23][13][17] <= img[10799];\
        in_img_array[23][14][0] <= img[10800];\
        in_img_array[23][14][1] <= img[10801];\
        in_img_array[23][14][2] <= img[10802];\
        in_img_array[23][14][3] <= img[10803];\
        in_img_array[23][14][4] <= img[10804];\
        in_img_array[23][14][5] <= img[10805];\
        in_img_array[23][14][6] <= img[10806];\
        in_img_array[23][14][7] <= img[10807];\
        in_img_array[23][14][8] <= img[10808];\
        in_img_array[23][14][9] <= img[10809];\
        in_img_array[23][14][10] <= img[10810];\
        in_img_array[23][14][11] <= img[10811];\
        in_img_array[23][14][12] <= img[10812];\
        in_img_array[23][14][13] <= img[10813];\
        in_img_array[23][14][14] <= img[10814];\
        in_img_array[23][14][15] <= img[10815];\
        in_img_array[23][14][16] <= img[10816];\
        in_img_array[23][14][17] <= img[10817];\
        in_img_array[23][15][0] <= img[10818];\
        in_img_array[23][15][1] <= img[10819];\
        in_img_array[23][15][2] <= img[10820];\
        in_img_array[23][15][3] <= img[10821];\
        in_img_array[23][15][4] <= img[10822];\
        in_img_array[23][15][5] <= img[10823];\
        in_img_array[23][15][6] <= img[10824];\
        in_img_array[23][15][7] <= img[10825];\
        in_img_array[23][15][8] <= img[10826];\
        in_img_array[23][15][9] <= img[10827];\
        in_img_array[23][15][10] <= img[10828];\
        in_img_array[23][15][11] <= img[10829];\
        in_img_array[23][15][12] <= img[10830];\
        in_img_array[23][15][13] <= img[10831];\
        in_img_array[23][15][14] <= img[10832];\
        in_img_array[23][15][15] <= img[10833];\
        in_img_array[23][15][16] <= img[10834];\
        in_img_array[23][15][17] <= img[10835];\
        in_img_array[23][16][0] <= img[10836];\
        in_img_array[23][16][1] <= img[10837];\
        in_img_array[23][16][2] <= img[10838];\
        in_img_array[23][16][3] <= img[10839];\
        in_img_array[23][16][4] <= img[10840];\
        in_img_array[23][16][5] <= img[10841];\
        in_img_array[23][16][6] <= img[10842];\
        in_img_array[23][16][7] <= img[10843];\
        in_img_array[23][16][8] <= img[10844];\
        in_img_array[23][16][9] <= img[10845];\
        in_img_array[23][16][10] <= img[10846];\
        in_img_array[23][16][11] <= img[10847];\
        in_img_array[23][16][12] <= img[10848];\
        in_img_array[23][16][13] <= img[10849];\
        in_img_array[23][16][14] <= img[10850];\
        in_img_array[23][16][15] <= img[10851];\
        in_img_array[23][16][16] <= img[10852];\
        in_img_array[23][16][17] <= img[10853];\
        in_img_array[23][17][0] <= img[10854];\
        in_img_array[23][17][1] <= img[10855];\
        in_img_array[23][17][2] <= img[10856];\
        in_img_array[23][17][3] <= img[10857];\
        in_img_array[23][17][4] <= img[10858];\
        in_img_array[23][17][5] <= img[10859];\
        in_img_array[23][17][6] <= img[10860];\
        in_img_array[23][17][7] <= img[10861];\
        in_img_array[23][17][8] <= img[10862];\
        in_img_array[23][17][9] <= img[10863];\
        in_img_array[23][17][10] <= img[10864];\
        in_img_array[23][17][11] <= img[10865];\
        in_img_array[23][17][12] <= img[10866];\
        in_img_array[23][17][13] <= img[10867];\
        in_img_array[23][17][14] <= img[10868];\
        in_img_array[23][17][15] <= img[10869];\
        in_img_array[23][17][16] <= img[10870];\
        in_img_array[23][17][17] <= img[10871];\
        in_img_array[23][18][0] <= img[10872];\
        in_img_array[23][18][1] <= img[10873];\
        in_img_array[23][18][2] <= img[10874];\
        in_img_array[23][18][3] <= img[10875];\
        in_img_array[23][18][4] <= img[10876];\
        in_img_array[23][18][5] <= img[10877];\
        in_img_array[23][18][6] <= img[10878];\
        in_img_array[23][18][7] <= img[10879];\
        in_img_array[23][18][8] <= img[10880];\
        in_img_array[23][18][9] <= img[10881];\
        in_img_array[23][18][10] <= img[10882];\
        in_img_array[23][18][11] <= img[10883];\
        in_img_array[23][18][12] <= img[10884];\
        in_img_array[23][18][13] <= img[10885];\
        in_img_array[23][18][14] <= img[10886];\
        in_img_array[23][18][15] <= img[10887];\
        in_img_array[23][18][16] <= img[10888];\
        in_img_array[23][18][17] <= img[10889];\
        in_img_array[23][19][0] <= img[10890];\
        in_img_array[23][19][1] <= img[10891];\
        in_img_array[23][19][2] <= img[10892];\
        in_img_array[23][19][3] <= img[10893];\
        in_img_array[23][19][4] <= img[10894];\
        in_img_array[23][19][5] <= img[10895];\
        in_img_array[23][19][6] <= img[10896];\
        in_img_array[23][19][7] <= img[10897];\
        in_img_array[23][19][8] <= img[10898];\
        in_img_array[23][19][9] <= img[10899];\
        in_img_array[23][19][10] <= img[10900];\
        in_img_array[23][19][11] <= img[10901];\
        in_img_array[23][19][12] <= img[10902];\
        in_img_array[23][19][13] <= img[10903];\
        in_img_array[23][19][14] <= img[10904];\
        in_img_array[23][19][15] <= img[10905];\
        in_img_array[23][19][16] <= img[10906];\
        in_img_array[23][19][17] <= img[10907];\
        in_img_array[23][20][0] <= img[10908];\
        in_img_array[23][20][1] <= img[10909];\
        in_img_array[23][20][2] <= img[10910];\
        in_img_array[23][20][3] <= img[10911];\
        in_img_array[23][20][4] <= img[10912];\
        in_img_array[23][20][5] <= img[10913];\
        in_img_array[23][20][6] <= img[10914];\
        in_img_array[23][20][7] <= img[10915];\
        in_img_array[23][20][8] <= img[10916];\
        in_img_array[23][20][9] <= img[10917];\
        in_img_array[23][20][10] <= img[10918];\
        in_img_array[23][20][11] <= img[10919];\
        in_img_array[23][20][12] <= img[10920];\
        in_img_array[23][20][13] <= img[10921];\
        in_img_array[23][20][14] <= img[10922];\
        in_img_array[23][20][15] <= img[10923];\
        in_img_array[23][20][16] <= img[10924];\
        in_img_array[23][20][17] <= img[10925];\
        in_img_array[23][21][0] <= img[10926];\
        in_img_array[23][21][1] <= img[10927];\
        in_img_array[23][21][2] <= img[10928];\
        in_img_array[23][21][3] <= img[10929];\
        in_img_array[23][21][4] <= img[10930];\
        in_img_array[23][21][5] <= img[10931];\
        in_img_array[23][21][6] <= img[10932];\
        in_img_array[23][21][7] <= img[10933];\
        in_img_array[23][21][8] <= img[10934];\
        in_img_array[23][21][9] <= img[10935];\
        in_img_array[23][21][10] <= img[10936];\
        in_img_array[23][21][11] <= img[10937];\
        in_img_array[23][21][12] <= img[10938];\
        in_img_array[23][21][13] <= img[10939];\
        in_img_array[23][21][14] <= img[10940];\
        in_img_array[23][21][15] <= img[10941];\
        in_img_array[23][21][16] <= img[10942];\
        in_img_array[23][21][17] <= img[10943];\
        in_img_array[23][22][0] <= img[10944];\
        in_img_array[23][22][1] <= img[10945];\
        in_img_array[23][22][2] <= img[10946];\
        in_img_array[23][22][3] <= img[10947];\
        in_img_array[23][22][4] <= img[10948];\
        in_img_array[23][22][5] <= img[10949];\
        in_img_array[23][22][6] <= img[10950];\
        in_img_array[23][22][7] <= img[10951];\
        in_img_array[23][22][8] <= img[10952];\
        in_img_array[23][22][9] <= img[10953];\
        in_img_array[23][22][10] <= img[10954];\
        in_img_array[23][22][11] <= img[10955];\
        in_img_array[23][22][12] <= img[10956];\
        in_img_array[23][22][13] <= img[10957];\
        in_img_array[23][22][14] <= img[10958];\
        in_img_array[23][22][15] <= img[10959];\
        in_img_array[23][22][16] <= img[10960];\
        in_img_array[23][22][17] <= img[10961];\
        in_img_array[23][23][0] <= img[10962];\
        in_img_array[23][23][1] <= img[10963];\
        in_img_array[23][23][2] <= img[10964];\
        in_img_array[23][23][3] <= img[10965];\
        in_img_array[23][23][4] <= img[10966];\
        in_img_array[23][23][5] <= img[10967];\
        in_img_array[23][23][6] <= img[10968];\
        in_img_array[23][23][7] <= img[10969];\
        in_img_array[23][23][8] <= img[10970];\
        in_img_array[23][23][9] <= img[10971];\
        in_img_array[23][23][10] <= img[10972];\
        in_img_array[23][23][11] <= img[10973];\
        in_img_array[23][23][12] <= img[10974];\
        in_img_array[23][23][13] <= img[10975];\
        in_img_array[23][23][14] <= img[10976];\
        in_img_array[23][23][15] <= img[10977];\
        in_img_array[23][23][16] <= img[10978];\
        in_img_array[23][23][17] <= img[10979];\
        in_img_array[23][24][0] <= img[10980];\
        in_img_array[23][24][1] <= img[10981];\
        in_img_array[23][24][2] <= img[10982];\
        in_img_array[23][24][3] <= img[10983];\
        in_img_array[23][24][4] <= img[10984];\
        in_img_array[23][24][5] <= img[10985];\
        in_img_array[23][24][6] <= img[10986];\
        in_img_array[23][24][7] <= img[10987];\
        in_img_array[23][24][8] <= img[10988];\
        in_img_array[23][24][9] <= img[10989];\
        in_img_array[23][24][10] <= img[10990];\
        in_img_array[23][24][11] <= img[10991];\
        in_img_array[23][24][12] <= img[10992];\
        in_img_array[23][24][13] <= img[10993];\
        in_img_array[23][24][14] <= img[10994];\
        in_img_array[23][24][15] <= img[10995];\
        in_img_array[23][24][16] <= img[10996];\
        in_img_array[23][24][17] <= img[10997];\
        in_img_array[23][25][0] <= img[10998];\
        in_img_array[23][25][1] <= img[10999];\
        in_img_array[23][25][2] <= img[11000];\
        in_img_array[23][25][3] <= img[11001];\
        in_img_array[23][25][4] <= img[11002];\
        in_img_array[23][25][5] <= img[11003];\
        in_img_array[23][25][6] <= img[11004];\
        in_img_array[23][25][7] <= img[11005];\
        in_img_array[23][25][8] <= img[11006];\
        in_img_array[23][25][9] <= img[11007];\
        in_img_array[23][25][10] <= img[11008];\
        in_img_array[23][25][11] <= img[11009];\
        in_img_array[23][25][12] <= img[11010];\
        in_img_array[23][25][13] <= img[11011];\
        in_img_array[23][25][14] <= img[11012];\
        in_img_array[23][25][15] <= img[11013];\
        in_img_array[23][25][16] <= img[11014];\
        in_img_array[23][25][17] <= img[11015];\
        in_img_array[23][26][0] <= img[11016];\
        in_img_array[23][26][1] <= img[11017];\
        in_img_array[23][26][2] <= img[11018];\
        in_img_array[23][26][3] <= img[11019];\
        in_img_array[23][26][4] <= img[11020];\
        in_img_array[23][26][5] <= img[11021];\
        in_img_array[23][26][6] <= img[11022];\
        in_img_array[23][26][7] <= img[11023];\
        in_img_array[23][26][8] <= img[11024];\
        in_img_array[23][26][9] <= img[11025];\
        in_img_array[23][26][10] <= img[11026];\
        in_img_array[23][26][11] <= img[11027];\
        in_img_array[23][26][12] <= img[11028];\
        in_img_array[23][26][13] <= img[11029];\
        in_img_array[23][26][14] <= img[11030];\
        in_img_array[23][26][15] <= img[11031];\
        in_img_array[23][26][16] <= img[11032];\
        in_img_array[23][26][17] <= img[11033];\
        in_img_array[23][27][0] <= img[11034];\
        in_img_array[23][27][1] <= img[11035];\
        in_img_array[23][27][2] <= img[11036];\
        in_img_array[23][27][3] <= img[11037];\
        in_img_array[23][27][4] <= img[11038];\
        in_img_array[23][27][5] <= img[11039];\
        in_img_array[23][27][6] <= img[11040];\
        in_img_array[23][27][7] <= img[11041];\
        in_img_array[23][27][8] <= img[11042];\
        in_img_array[23][27][9] <= img[11043];\
        in_img_array[23][27][10] <= img[11044];\
        in_img_array[23][27][11] <= img[11045];\
        in_img_array[23][27][12] <= img[11046];\
        in_img_array[23][27][13] <= img[11047];\
        in_img_array[23][27][14] <= img[11048];\
        in_img_array[23][27][15] <= img[11049];\
        in_img_array[23][27][16] <= img[11050];\
        in_img_array[23][27][17] <= img[11051];\
        in_img_array[23][28][0] <= img[11052];\
        in_img_array[23][28][1] <= img[11053];\
        in_img_array[23][28][2] <= img[11054];\
        in_img_array[23][28][3] <= img[11055];\
        in_img_array[23][28][4] <= img[11056];\
        in_img_array[23][28][5] <= img[11057];\
        in_img_array[23][28][6] <= img[11058];\
        in_img_array[23][28][7] <= img[11059];\
        in_img_array[23][28][8] <= img[11060];\
        in_img_array[23][28][9] <= img[11061];\
        in_img_array[23][28][10] <= img[11062];\
        in_img_array[23][28][11] <= img[11063];\
        in_img_array[23][28][12] <= img[11064];\
        in_img_array[23][28][13] <= img[11065];\
        in_img_array[23][28][14] <= img[11066];\
        in_img_array[23][28][15] <= img[11067];\
        in_img_array[23][28][16] <= img[11068];\
        in_img_array[23][28][17] <= img[11069];\
        in_img_array[23][29][0] <= img[11070];\
        in_img_array[23][29][1] <= img[11071];\
        in_img_array[23][29][2] <= img[11072];\
        in_img_array[23][29][3] <= img[11073];\
        in_img_array[23][29][4] <= img[11074];\
        in_img_array[23][29][5] <= img[11075];\
        in_img_array[23][29][6] <= img[11076];\
        in_img_array[23][29][7] <= img[11077];\
        in_img_array[23][29][8] <= img[11078];\
        in_img_array[23][29][9] <= img[11079];\
        in_img_array[23][29][10] <= img[11080];\
        in_img_array[23][29][11] <= img[11081];\
        in_img_array[23][29][12] <= img[11082];\
        in_img_array[23][29][13] <= img[11083];\
        in_img_array[23][29][14] <= img[11084];\
        in_img_array[23][29][15] <= img[11085];\
        in_img_array[23][29][16] <= img[11086];\
        in_img_array[23][29][17] <= img[11087];\
        in_img_array[24][2][0] <= img[11088];\
        in_img_array[24][2][1] <= img[11089];\
        in_img_array[24][2][2] <= img[11090];\
        in_img_array[24][2][3] <= img[11091];\
        in_img_array[24][2][4] <= img[11092];\
        in_img_array[24][2][5] <= img[11093];\
        in_img_array[24][2][6] <= img[11094];\
        in_img_array[24][2][7] <= img[11095];\
        in_img_array[24][2][8] <= img[11096];\
        in_img_array[24][2][9] <= img[11097];\
        in_img_array[24][2][10] <= img[11098];\
        in_img_array[24][2][11] <= img[11099];\
        in_img_array[24][2][12] <= img[11100];\
        in_img_array[24][2][13] <= img[11101];\
        in_img_array[24][2][14] <= img[11102];\
        in_img_array[24][2][15] <= img[11103];\
        in_img_array[24][2][16] <= img[11104];\
        in_img_array[24][2][17] <= img[11105];\
        in_img_array[24][3][0] <= img[11106];\
        in_img_array[24][3][1] <= img[11107];\
        in_img_array[24][3][2] <= img[11108];\
        in_img_array[24][3][3] <= img[11109];\
        in_img_array[24][3][4] <= img[11110];\
        in_img_array[24][3][5] <= img[11111];\
        in_img_array[24][3][6] <= img[11112];\
        in_img_array[24][3][7] <= img[11113];\
        in_img_array[24][3][8] <= img[11114];\
        in_img_array[24][3][9] <= img[11115];\
        in_img_array[24][3][10] <= img[11116];\
        in_img_array[24][3][11] <= img[11117];\
        in_img_array[24][3][12] <= img[11118];\
        in_img_array[24][3][13] <= img[11119];\
        in_img_array[24][3][14] <= img[11120];\
        in_img_array[24][3][15] <= img[11121];\
        in_img_array[24][3][16] <= img[11122];\
        in_img_array[24][3][17] <= img[11123];\
        in_img_array[24][4][0] <= img[11124];\
        in_img_array[24][4][1] <= img[11125];\
        in_img_array[24][4][2] <= img[11126];\
        in_img_array[24][4][3] <= img[11127];\
        in_img_array[24][4][4] <= img[11128];\
        in_img_array[24][4][5] <= img[11129];\
        in_img_array[24][4][6] <= img[11130];\
        in_img_array[24][4][7] <= img[11131];\
        in_img_array[24][4][8] <= img[11132];\
        in_img_array[24][4][9] <= img[11133];\
        in_img_array[24][4][10] <= img[11134];\
        in_img_array[24][4][11] <= img[11135];\
        in_img_array[24][4][12] <= img[11136];\
        in_img_array[24][4][13] <= img[11137];\
        in_img_array[24][4][14] <= img[11138];\
        in_img_array[24][4][15] <= img[11139];\
        in_img_array[24][4][16] <= img[11140];\
        in_img_array[24][4][17] <= img[11141];\
        in_img_array[24][5][0] <= img[11142];\
        in_img_array[24][5][1] <= img[11143];\
        in_img_array[24][5][2] <= img[11144];\
        in_img_array[24][5][3] <= img[11145];\
        in_img_array[24][5][4] <= img[11146];\
        in_img_array[24][5][5] <= img[11147];\
        in_img_array[24][5][6] <= img[11148];\
        in_img_array[24][5][7] <= img[11149];\
        in_img_array[24][5][8] <= img[11150];\
        in_img_array[24][5][9] <= img[11151];\
        in_img_array[24][5][10] <= img[11152];\
        in_img_array[24][5][11] <= img[11153];\
        in_img_array[24][5][12] <= img[11154];\
        in_img_array[24][5][13] <= img[11155];\
        in_img_array[24][5][14] <= img[11156];\
        in_img_array[24][5][15] <= img[11157];\
        in_img_array[24][5][16] <= img[11158];\
        in_img_array[24][5][17] <= img[11159];\
        in_img_array[24][6][0] <= img[11160];\
        in_img_array[24][6][1] <= img[11161];\
        in_img_array[24][6][2] <= img[11162];\
        in_img_array[24][6][3] <= img[11163];\
        in_img_array[24][6][4] <= img[11164];\
        in_img_array[24][6][5] <= img[11165];\
        in_img_array[24][6][6] <= img[11166];\
        in_img_array[24][6][7] <= img[11167];\
        in_img_array[24][6][8] <= img[11168];\
        in_img_array[24][6][9] <= img[11169];\
        in_img_array[24][6][10] <= img[11170];\
        in_img_array[24][6][11] <= img[11171];\
        in_img_array[24][6][12] <= img[11172];\
        in_img_array[24][6][13] <= img[11173];\
        in_img_array[24][6][14] <= img[11174];\
        in_img_array[24][6][15] <= img[11175];\
        in_img_array[24][6][16] <= img[11176];\
        in_img_array[24][6][17] <= img[11177];\
        in_img_array[24][7][0] <= img[11178];\
        in_img_array[24][7][1] <= img[11179];\
        in_img_array[24][7][2] <= img[11180];\
        in_img_array[24][7][3] <= img[11181];\
        in_img_array[24][7][4] <= img[11182];\
        in_img_array[24][7][5] <= img[11183];\
        in_img_array[24][7][6] <= img[11184];\
        in_img_array[24][7][7] <= img[11185];\
        in_img_array[24][7][8] <= img[11186];\
        in_img_array[24][7][9] <= img[11187];\
        in_img_array[24][7][10] <= img[11188];\
        in_img_array[24][7][11] <= img[11189];\
        in_img_array[24][7][12] <= img[11190];\
        in_img_array[24][7][13] <= img[11191];\
        in_img_array[24][7][14] <= img[11192];\
        in_img_array[24][7][15] <= img[11193];\
        in_img_array[24][7][16] <= img[11194];\
        in_img_array[24][7][17] <= img[11195];\
        in_img_array[24][8][0] <= img[11196];\
        in_img_array[24][8][1] <= img[11197];\
        in_img_array[24][8][2] <= img[11198];\
        in_img_array[24][8][3] <= img[11199];\
        in_img_array[24][8][4] <= img[11200];\
        in_img_array[24][8][5] <= img[11201];\
        in_img_array[24][8][6] <= img[11202];\
        in_img_array[24][8][7] <= img[11203];\
        in_img_array[24][8][8] <= img[11204];\
        in_img_array[24][8][9] <= img[11205];\
        in_img_array[24][8][10] <= img[11206];\
        in_img_array[24][8][11] <= img[11207];\
        in_img_array[24][8][12] <= img[11208];\
        in_img_array[24][8][13] <= img[11209];\
        in_img_array[24][8][14] <= img[11210];\
        in_img_array[24][8][15] <= img[11211];\
        in_img_array[24][8][16] <= img[11212];\
        in_img_array[24][8][17] <= img[11213];\
        in_img_array[24][9][0] <= img[11214];\
        in_img_array[24][9][1] <= img[11215];\
        in_img_array[24][9][2] <= img[11216];\
        in_img_array[24][9][3] <= img[11217];\
        in_img_array[24][9][4] <= img[11218];\
        in_img_array[24][9][5] <= img[11219];\
        in_img_array[24][9][6] <= img[11220];\
        in_img_array[24][9][7] <= img[11221];\
        in_img_array[24][9][8] <= img[11222];\
        in_img_array[24][9][9] <= img[11223];\
        in_img_array[24][9][10] <= img[11224];\
        in_img_array[24][9][11] <= img[11225];\
        in_img_array[24][9][12] <= img[11226];\
        in_img_array[24][9][13] <= img[11227];\
        in_img_array[24][9][14] <= img[11228];\
        in_img_array[24][9][15] <= img[11229];\
        in_img_array[24][9][16] <= img[11230];\
        in_img_array[24][9][17] <= img[11231];\
        in_img_array[24][10][0] <= img[11232];\
        in_img_array[24][10][1] <= img[11233];\
        in_img_array[24][10][2] <= img[11234];\
        in_img_array[24][10][3] <= img[11235];\
        in_img_array[24][10][4] <= img[11236];\
        in_img_array[24][10][5] <= img[11237];\
        in_img_array[24][10][6] <= img[11238];\
        in_img_array[24][10][7] <= img[11239];\
        in_img_array[24][10][8] <= img[11240];\
        in_img_array[24][10][9] <= img[11241];\
        in_img_array[24][10][10] <= img[11242];\
        in_img_array[24][10][11] <= img[11243];\
        in_img_array[24][10][12] <= img[11244];\
        in_img_array[24][10][13] <= img[11245];\
        in_img_array[24][10][14] <= img[11246];\
        in_img_array[24][10][15] <= img[11247];\
        in_img_array[24][10][16] <= img[11248];\
        in_img_array[24][10][17] <= img[11249];\
        in_img_array[24][11][0] <= img[11250];\
        in_img_array[24][11][1] <= img[11251];\
        in_img_array[24][11][2] <= img[11252];\
        in_img_array[24][11][3] <= img[11253];\
        in_img_array[24][11][4] <= img[11254];\
        in_img_array[24][11][5] <= img[11255];\
        in_img_array[24][11][6] <= img[11256];\
        in_img_array[24][11][7] <= img[11257];\
        in_img_array[24][11][8] <= img[11258];\
        in_img_array[24][11][9] <= img[11259];\
        in_img_array[24][11][10] <= img[11260];\
        in_img_array[24][11][11] <= img[11261];\
        in_img_array[24][11][12] <= img[11262];\
        in_img_array[24][11][13] <= img[11263];\
        in_img_array[24][11][14] <= img[11264];\
        in_img_array[24][11][15] <= img[11265];\
        in_img_array[24][11][16] <= img[11266];\
        in_img_array[24][11][17] <= img[11267];\
        in_img_array[24][12][0] <= img[11268];\
        in_img_array[24][12][1] <= img[11269];\
        in_img_array[24][12][2] <= img[11270];\
        in_img_array[24][12][3] <= img[11271];\
        in_img_array[24][12][4] <= img[11272];\
        in_img_array[24][12][5] <= img[11273];\
        in_img_array[24][12][6] <= img[11274];\
        in_img_array[24][12][7] <= img[11275];\
        in_img_array[24][12][8] <= img[11276];\
        in_img_array[24][12][9] <= img[11277];\
        in_img_array[24][12][10] <= img[11278];\
        in_img_array[24][12][11] <= img[11279];\
        in_img_array[24][12][12] <= img[11280];\
        in_img_array[24][12][13] <= img[11281];\
        in_img_array[24][12][14] <= img[11282];\
        in_img_array[24][12][15] <= img[11283];\
        in_img_array[24][12][16] <= img[11284];\
        in_img_array[24][12][17] <= img[11285];\
        in_img_array[24][13][0] <= img[11286];\
        in_img_array[24][13][1] <= img[11287];\
        in_img_array[24][13][2] <= img[11288];\
        in_img_array[24][13][3] <= img[11289];\
        in_img_array[24][13][4] <= img[11290];\
        in_img_array[24][13][5] <= img[11291];\
        in_img_array[24][13][6] <= img[11292];\
        in_img_array[24][13][7] <= img[11293];\
        in_img_array[24][13][8] <= img[11294];\
        in_img_array[24][13][9] <= img[11295];\
        in_img_array[24][13][10] <= img[11296];\
        in_img_array[24][13][11] <= img[11297];\
        in_img_array[24][13][12] <= img[11298];\
        in_img_array[24][13][13] <= img[11299];\
        in_img_array[24][13][14] <= img[11300];\
        in_img_array[24][13][15] <= img[11301];\
        in_img_array[24][13][16] <= img[11302];\
        in_img_array[24][13][17] <= img[11303];\
        in_img_array[24][14][0] <= img[11304];\
        in_img_array[24][14][1] <= img[11305];\
        in_img_array[24][14][2] <= img[11306];\
        in_img_array[24][14][3] <= img[11307];\
        in_img_array[24][14][4] <= img[11308];\
        in_img_array[24][14][5] <= img[11309];\
        in_img_array[24][14][6] <= img[11310];\
        in_img_array[24][14][7] <= img[11311];\
        in_img_array[24][14][8] <= img[11312];\
        in_img_array[24][14][9] <= img[11313];\
        in_img_array[24][14][10] <= img[11314];\
        in_img_array[24][14][11] <= img[11315];\
        in_img_array[24][14][12] <= img[11316];\
        in_img_array[24][14][13] <= img[11317];\
        in_img_array[24][14][14] <= img[11318];\
        in_img_array[24][14][15] <= img[11319];\
        in_img_array[24][14][16] <= img[11320];\
        in_img_array[24][14][17] <= img[11321];\
        in_img_array[24][15][0] <= img[11322];\
        in_img_array[24][15][1] <= img[11323];\
        in_img_array[24][15][2] <= img[11324];\
        in_img_array[24][15][3] <= img[11325];\
        in_img_array[24][15][4] <= img[11326];\
        in_img_array[24][15][5] <= img[11327];\
        in_img_array[24][15][6] <= img[11328];\
        in_img_array[24][15][7] <= img[11329];\
        in_img_array[24][15][8] <= img[11330];\
        in_img_array[24][15][9] <= img[11331];\
        in_img_array[24][15][10] <= img[11332];\
        in_img_array[24][15][11] <= img[11333];\
        in_img_array[24][15][12] <= img[11334];\
        in_img_array[24][15][13] <= img[11335];\
        in_img_array[24][15][14] <= img[11336];\
        in_img_array[24][15][15] <= img[11337];\
        in_img_array[24][15][16] <= img[11338];\
        in_img_array[24][15][17] <= img[11339];\
        in_img_array[24][16][0] <= img[11340];\
        in_img_array[24][16][1] <= img[11341];\
        in_img_array[24][16][2] <= img[11342];\
        in_img_array[24][16][3] <= img[11343];\
        in_img_array[24][16][4] <= img[11344];\
        in_img_array[24][16][5] <= img[11345];\
        in_img_array[24][16][6] <= img[11346];\
        in_img_array[24][16][7] <= img[11347];\
        in_img_array[24][16][8] <= img[11348];\
        in_img_array[24][16][9] <= img[11349];\
        in_img_array[24][16][10] <= img[11350];\
        in_img_array[24][16][11] <= img[11351];\
        in_img_array[24][16][12] <= img[11352];\
        in_img_array[24][16][13] <= img[11353];\
        in_img_array[24][16][14] <= img[11354];\
        in_img_array[24][16][15] <= img[11355];\
        in_img_array[24][16][16] <= img[11356];\
        in_img_array[24][16][17] <= img[11357];\
        in_img_array[24][17][0] <= img[11358];\
        in_img_array[24][17][1] <= img[11359];\
        in_img_array[24][17][2] <= img[11360];\
        in_img_array[24][17][3] <= img[11361];\
        in_img_array[24][17][4] <= img[11362];\
        in_img_array[24][17][5] <= img[11363];\
        in_img_array[24][17][6] <= img[11364];\
        in_img_array[24][17][7] <= img[11365];\
        in_img_array[24][17][8] <= img[11366];\
        in_img_array[24][17][9] <= img[11367];\
        in_img_array[24][17][10] <= img[11368];\
        in_img_array[24][17][11] <= img[11369];\
        in_img_array[24][17][12] <= img[11370];\
        in_img_array[24][17][13] <= img[11371];\
        in_img_array[24][17][14] <= img[11372];\
        in_img_array[24][17][15] <= img[11373];\
        in_img_array[24][17][16] <= img[11374];\
        in_img_array[24][17][17] <= img[11375];\
        in_img_array[24][18][0] <= img[11376];\
        in_img_array[24][18][1] <= img[11377];\
        in_img_array[24][18][2] <= img[11378];\
        in_img_array[24][18][3] <= img[11379];\
        in_img_array[24][18][4] <= img[11380];\
        in_img_array[24][18][5] <= img[11381];\
        in_img_array[24][18][6] <= img[11382];\
        in_img_array[24][18][7] <= img[11383];\
        in_img_array[24][18][8] <= img[11384];\
        in_img_array[24][18][9] <= img[11385];\
        in_img_array[24][18][10] <= img[11386];\
        in_img_array[24][18][11] <= img[11387];\
        in_img_array[24][18][12] <= img[11388];\
        in_img_array[24][18][13] <= img[11389];\
        in_img_array[24][18][14] <= img[11390];\
        in_img_array[24][18][15] <= img[11391];\
        in_img_array[24][18][16] <= img[11392];\
        in_img_array[24][18][17] <= img[11393];\
        in_img_array[24][19][0] <= img[11394];\
        in_img_array[24][19][1] <= img[11395];\
        in_img_array[24][19][2] <= img[11396];\
        in_img_array[24][19][3] <= img[11397];\
        in_img_array[24][19][4] <= img[11398];\
        in_img_array[24][19][5] <= img[11399];\
        in_img_array[24][19][6] <= img[11400];\
        in_img_array[24][19][7] <= img[11401];\
        in_img_array[24][19][8] <= img[11402];\
        in_img_array[24][19][9] <= img[11403];\
        in_img_array[24][19][10] <= img[11404];\
        in_img_array[24][19][11] <= img[11405];\
        in_img_array[24][19][12] <= img[11406];\
        in_img_array[24][19][13] <= img[11407];\
        in_img_array[24][19][14] <= img[11408];\
        in_img_array[24][19][15] <= img[11409];\
        in_img_array[24][19][16] <= img[11410];\
        in_img_array[24][19][17] <= img[11411];\
        in_img_array[24][20][0] <= img[11412];\
        in_img_array[24][20][1] <= img[11413];\
        in_img_array[24][20][2] <= img[11414];\
        in_img_array[24][20][3] <= img[11415];\
        in_img_array[24][20][4] <= img[11416];\
        in_img_array[24][20][5] <= img[11417];\
        in_img_array[24][20][6] <= img[11418];\
        in_img_array[24][20][7] <= img[11419];\
        in_img_array[24][20][8] <= img[11420];\
        in_img_array[24][20][9] <= img[11421];\
        in_img_array[24][20][10] <= img[11422];\
        in_img_array[24][20][11] <= img[11423];\
        in_img_array[24][20][12] <= img[11424];\
        in_img_array[24][20][13] <= img[11425];\
        in_img_array[24][20][14] <= img[11426];\
        in_img_array[24][20][15] <= img[11427];\
        in_img_array[24][20][16] <= img[11428];\
        in_img_array[24][20][17] <= img[11429];\
        in_img_array[24][21][0] <= img[11430];\
        in_img_array[24][21][1] <= img[11431];\
        in_img_array[24][21][2] <= img[11432];\
        in_img_array[24][21][3] <= img[11433];\
        in_img_array[24][21][4] <= img[11434];\
        in_img_array[24][21][5] <= img[11435];\
        in_img_array[24][21][6] <= img[11436];\
        in_img_array[24][21][7] <= img[11437];\
        in_img_array[24][21][8] <= img[11438];\
        in_img_array[24][21][9] <= img[11439];\
        in_img_array[24][21][10] <= img[11440];\
        in_img_array[24][21][11] <= img[11441];\
        in_img_array[24][21][12] <= img[11442];\
        in_img_array[24][21][13] <= img[11443];\
        in_img_array[24][21][14] <= img[11444];\
        in_img_array[24][21][15] <= img[11445];\
        in_img_array[24][21][16] <= img[11446];\
        in_img_array[24][21][17] <= img[11447];\
        in_img_array[24][22][0] <= img[11448];\
        in_img_array[24][22][1] <= img[11449];\
        in_img_array[24][22][2] <= img[11450];\
        in_img_array[24][22][3] <= img[11451];\
        in_img_array[24][22][4] <= img[11452];\
        in_img_array[24][22][5] <= img[11453];\
        in_img_array[24][22][6] <= img[11454];\
        in_img_array[24][22][7] <= img[11455];\
        in_img_array[24][22][8] <= img[11456];\
        in_img_array[24][22][9] <= img[11457];\
        in_img_array[24][22][10] <= img[11458];\
        in_img_array[24][22][11] <= img[11459];\
        in_img_array[24][22][12] <= img[11460];\
        in_img_array[24][22][13] <= img[11461];\
        in_img_array[24][22][14] <= img[11462];\
        in_img_array[24][22][15] <= img[11463];\
        in_img_array[24][22][16] <= img[11464];\
        in_img_array[24][22][17] <= img[11465];\
        in_img_array[24][23][0] <= img[11466];\
        in_img_array[24][23][1] <= img[11467];\
        in_img_array[24][23][2] <= img[11468];\
        in_img_array[24][23][3] <= img[11469];\
        in_img_array[24][23][4] <= img[11470];\
        in_img_array[24][23][5] <= img[11471];\
        in_img_array[24][23][6] <= img[11472];\
        in_img_array[24][23][7] <= img[11473];\
        in_img_array[24][23][8] <= img[11474];\
        in_img_array[24][23][9] <= img[11475];\
        in_img_array[24][23][10] <= img[11476];\
        in_img_array[24][23][11] <= img[11477];\
        in_img_array[24][23][12] <= img[11478];\
        in_img_array[24][23][13] <= img[11479];\
        in_img_array[24][23][14] <= img[11480];\
        in_img_array[24][23][15] <= img[11481];\
        in_img_array[24][23][16] <= img[11482];\
        in_img_array[24][23][17] <= img[11483];\
        in_img_array[24][24][0] <= img[11484];\
        in_img_array[24][24][1] <= img[11485];\
        in_img_array[24][24][2] <= img[11486];\
        in_img_array[24][24][3] <= img[11487];\
        in_img_array[24][24][4] <= img[11488];\
        in_img_array[24][24][5] <= img[11489];\
        in_img_array[24][24][6] <= img[11490];\
        in_img_array[24][24][7] <= img[11491];\
        in_img_array[24][24][8] <= img[11492];\
        in_img_array[24][24][9] <= img[11493];\
        in_img_array[24][24][10] <= img[11494];\
        in_img_array[24][24][11] <= img[11495];\
        in_img_array[24][24][12] <= img[11496];\
        in_img_array[24][24][13] <= img[11497];\
        in_img_array[24][24][14] <= img[11498];\
        in_img_array[24][24][15] <= img[11499];\
        in_img_array[24][24][16] <= img[11500];\
        in_img_array[24][24][17] <= img[11501];\
        in_img_array[24][25][0] <= img[11502];\
        in_img_array[24][25][1] <= img[11503];\
        in_img_array[24][25][2] <= img[11504];\
        in_img_array[24][25][3] <= img[11505];\
        in_img_array[24][25][4] <= img[11506];\
        in_img_array[24][25][5] <= img[11507];\
        in_img_array[24][25][6] <= img[11508];\
        in_img_array[24][25][7] <= img[11509];\
        in_img_array[24][25][8] <= img[11510];\
        in_img_array[24][25][9] <= img[11511];\
        in_img_array[24][25][10] <= img[11512];\
        in_img_array[24][25][11] <= img[11513];\
        in_img_array[24][25][12] <= img[11514];\
        in_img_array[24][25][13] <= img[11515];\
        in_img_array[24][25][14] <= img[11516];\
        in_img_array[24][25][15] <= img[11517];\
        in_img_array[24][25][16] <= img[11518];\
        in_img_array[24][25][17] <= img[11519];\
        in_img_array[24][26][0] <= img[11520];\
        in_img_array[24][26][1] <= img[11521];\
        in_img_array[24][26][2] <= img[11522];\
        in_img_array[24][26][3] <= img[11523];\
        in_img_array[24][26][4] <= img[11524];\
        in_img_array[24][26][5] <= img[11525];\
        in_img_array[24][26][6] <= img[11526];\
        in_img_array[24][26][7] <= img[11527];\
        in_img_array[24][26][8] <= img[11528];\
        in_img_array[24][26][9] <= img[11529];\
        in_img_array[24][26][10] <= img[11530];\
        in_img_array[24][26][11] <= img[11531];\
        in_img_array[24][26][12] <= img[11532];\
        in_img_array[24][26][13] <= img[11533];\
        in_img_array[24][26][14] <= img[11534];\
        in_img_array[24][26][15] <= img[11535];\
        in_img_array[24][26][16] <= img[11536];\
        in_img_array[24][26][17] <= img[11537];\
        in_img_array[24][27][0] <= img[11538];\
        in_img_array[24][27][1] <= img[11539];\
        in_img_array[24][27][2] <= img[11540];\
        in_img_array[24][27][3] <= img[11541];\
        in_img_array[24][27][4] <= img[11542];\
        in_img_array[24][27][5] <= img[11543];\
        in_img_array[24][27][6] <= img[11544];\
        in_img_array[24][27][7] <= img[11545];\
        in_img_array[24][27][8] <= img[11546];\
        in_img_array[24][27][9] <= img[11547];\
        in_img_array[24][27][10] <= img[11548];\
        in_img_array[24][27][11] <= img[11549];\
        in_img_array[24][27][12] <= img[11550];\
        in_img_array[24][27][13] <= img[11551];\
        in_img_array[24][27][14] <= img[11552];\
        in_img_array[24][27][15] <= img[11553];\
        in_img_array[24][27][16] <= img[11554];\
        in_img_array[24][27][17] <= img[11555];\
        in_img_array[24][28][0] <= img[11556];\
        in_img_array[24][28][1] <= img[11557];\
        in_img_array[24][28][2] <= img[11558];\
        in_img_array[24][28][3] <= img[11559];\
        in_img_array[24][28][4] <= img[11560];\
        in_img_array[24][28][5] <= img[11561];\
        in_img_array[24][28][6] <= img[11562];\
        in_img_array[24][28][7] <= img[11563];\
        in_img_array[24][28][8] <= img[11564];\
        in_img_array[24][28][9] <= img[11565];\
        in_img_array[24][28][10] <= img[11566];\
        in_img_array[24][28][11] <= img[11567];\
        in_img_array[24][28][12] <= img[11568];\
        in_img_array[24][28][13] <= img[11569];\
        in_img_array[24][28][14] <= img[11570];\
        in_img_array[24][28][15] <= img[11571];\
        in_img_array[24][28][16] <= img[11572];\
        in_img_array[24][28][17] <= img[11573];\
        in_img_array[24][29][0] <= img[11574];\
        in_img_array[24][29][1] <= img[11575];\
        in_img_array[24][29][2] <= img[11576];\
        in_img_array[24][29][3] <= img[11577];\
        in_img_array[24][29][4] <= img[11578];\
        in_img_array[24][29][5] <= img[11579];\
        in_img_array[24][29][6] <= img[11580];\
        in_img_array[24][29][7] <= img[11581];\
        in_img_array[24][29][8] <= img[11582];\
        in_img_array[24][29][9] <= img[11583];\
        in_img_array[24][29][10] <= img[11584];\
        in_img_array[24][29][11] <= img[11585];\
        in_img_array[24][29][12] <= img[11586];\
        in_img_array[24][29][13] <= img[11587];\
        in_img_array[24][29][14] <= img[11588];\
        in_img_array[24][29][15] <= img[11589];\
        in_img_array[24][29][16] <= img[11590];\
        in_img_array[24][29][17] <= img[11591];\
        in_img_array[25][2][0] <= img[11592];\
        in_img_array[25][2][1] <= img[11593];\
        in_img_array[25][2][2] <= img[11594];\
        in_img_array[25][2][3] <= img[11595];\
        in_img_array[25][2][4] <= img[11596];\
        in_img_array[25][2][5] <= img[11597];\
        in_img_array[25][2][6] <= img[11598];\
        in_img_array[25][2][7] <= img[11599];\
        in_img_array[25][2][8] <= img[11600];\
        in_img_array[25][2][9] <= img[11601];\
        in_img_array[25][2][10] <= img[11602];\
        in_img_array[25][2][11] <= img[11603];\
        in_img_array[25][2][12] <= img[11604];\
        in_img_array[25][2][13] <= img[11605];\
        in_img_array[25][2][14] <= img[11606];\
        in_img_array[25][2][15] <= img[11607];\
        in_img_array[25][2][16] <= img[11608];\
        in_img_array[25][2][17] <= img[11609];\
        in_img_array[25][3][0] <= img[11610];\
        in_img_array[25][3][1] <= img[11611];\
        in_img_array[25][3][2] <= img[11612];\
        in_img_array[25][3][3] <= img[11613];\
        in_img_array[25][3][4] <= img[11614];\
        in_img_array[25][3][5] <= img[11615];\
        in_img_array[25][3][6] <= img[11616];\
        in_img_array[25][3][7] <= img[11617];\
        in_img_array[25][3][8] <= img[11618];\
        in_img_array[25][3][9] <= img[11619];\
        in_img_array[25][3][10] <= img[11620];\
        in_img_array[25][3][11] <= img[11621];\
        in_img_array[25][3][12] <= img[11622];\
        in_img_array[25][3][13] <= img[11623];\
        in_img_array[25][3][14] <= img[11624];\
        in_img_array[25][3][15] <= img[11625];\
        in_img_array[25][3][16] <= img[11626];\
        in_img_array[25][3][17] <= img[11627];\
        in_img_array[25][4][0] <= img[11628];\
        in_img_array[25][4][1] <= img[11629];\
        in_img_array[25][4][2] <= img[11630];\
        in_img_array[25][4][3] <= img[11631];\
        in_img_array[25][4][4] <= img[11632];\
        in_img_array[25][4][5] <= img[11633];\
        in_img_array[25][4][6] <= img[11634];\
        in_img_array[25][4][7] <= img[11635];\
        in_img_array[25][4][8] <= img[11636];\
        in_img_array[25][4][9] <= img[11637];\
        in_img_array[25][4][10] <= img[11638];\
        in_img_array[25][4][11] <= img[11639];\
        in_img_array[25][4][12] <= img[11640];\
        in_img_array[25][4][13] <= img[11641];\
        in_img_array[25][4][14] <= img[11642];\
        in_img_array[25][4][15] <= img[11643];\
        in_img_array[25][4][16] <= img[11644];\
        in_img_array[25][4][17] <= img[11645];\
        in_img_array[25][5][0] <= img[11646];\
        in_img_array[25][5][1] <= img[11647];\
        in_img_array[25][5][2] <= img[11648];\
        in_img_array[25][5][3] <= img[11649];\
        in_img_array[25][5][4] <= img[11650];\
        in_img_array[25][5][5] <= img[11651];\
        in_img_array[25][5][6] <= img[11652];\
        in_img_array[25][5][7] <= img[11653];\
        in_img_array[25][5][8] <= img[11654];\
        in_img_array[25][5][9] <= img[11655];\
        in_img_array[25][5][10] <= img[11656];\
        in_img_array[25][5][11] <= img[11657];\
        in_img_array[25][5][12] <= img[11658];\
        in_img_array[25][5][13] <= img[11659];\
        in_img_array[25][5][14] <= img[11660];\
        in_img_array[25][5][15] <= img[11661];\
        in_img_array[25][5][16] <= img[11662];\
        in_img_array[25][5][17] <= img[11663];\
        in_img_array[25][6][0] <= img[11664];\
        in_img_array[25][6][1] <= img[11665];\
        in_img_array[25][6][2] <= img[11666];\
        in_img_array[25][6][3] <= img[11667];\
        in_img_array[25][6][4] <= img[11668];\
        in_img_array[25][6][5] <= img[11669];\
        in_img_array[25][6][6] <= img[11670];\
        in_img_array[25][6][7] <= img[11671];\
        in_img_array[25][6][8] <= img[11672];\
        in_img_array[25][6][9] <= img[11673];\
        in_img_array[25][6][10] <= img[11674];\
        in_img_array[25][6][11] <= img[11675];\
        in_img_array[25][6][12] <= img[11676];\
        in_img_array[25][6][13] <= img[11677];\
        in_img_array[25][6][14] <= img[11678];\
        in_img_array[25][6][15] <= img[11679];\
        in_img_array[25][6][16] <= img[11680];\
        in_img_array[25][6][17] <= img[11681];\
        in_img_array[25][7][0] <= img[11682];\
        in_img_array[25][7][1] <= img[11683];\
        in_img_array[25][7][2] <= img[11684];\
        in_img_array[25][7][3] <= img[11685];\
        in_img_array[25][7][4] <= img[11686];\
        in_img_array[25][7][5] <= img[11687];\
        in_img_array[25][7][6] <= img[11688];\
        in_img_array[25][7][7] <= img[11689];\
        in_img_array[25][7][8] <= img[11690];\
        in_img_array[25][7][9] <= img[11691];\
        in_img_array[25][7][10] <= img[11692];\
        in_img_array[25][7][11] <= img[11693];\
        in_img_array[25][7][12] <= img[11694];\
        in_img_array[25][7][13] <= img[11695];\
        in_img_array[25][7][14] <= img[11696];\
        in_img_array[25][7][15] <= img[11697];\
        in_img_array[25][7][16] <= img[11698];\
        in_img_array[25][7][17] <= img[11699];\
        in_img_array[25][8][0] <= img[11700];\
        in_img_array[25][8][1] <= img[11701];\
        in_img_array[25][8][2] <= img[11702];\
        in_img_array[25][8][3] <= img[11703];\
        in_img_array[25][8][4] <= img[11704];\
        in_img_array[25][8][5] <= img[11705];\
        in_img_array[25][8][6] <= img[11706];\
        in_img_array[25][8][7] <= img[11707];\
        in_img_array[25][8][8] <= img[11708];\
        in_img_array[25][8][9] <= img[11709];\
        in_img_array[25][8][10] <= img[11710];\
        in_img_array[25][8][11] <= img[11711];\
        in_img_array[25][8][12] <= img[11712];\
        in_img_array[25][8][13] <= img[11713];\
        in_img_array[25][8][14] <= img[11714];\
        in_img_array[25][8][15] <= img[11715];\
        in_img_array[25][8][16] <= img[11716];\
        in_img_array[25][8][17] <= img[11717];\
        in_img_array[25][9][0] <= img[11718];\
        in_img_array[25][9][1] <= img[11719];\
        in_img_array[25][9][2] <= img[11720];\
        in_img_array[25][9][3] <= img[11721];\
        in_img_array[25][9][4] <= img[11722];\
        in_img_array[25][9][5] <= img[11723];\
        in_img_array[25][9][6] <= img[11724];\
        in_img_array[25][9][7] <= img[11725];\
        in_img_array[25][9][8] <= img[11726];\
        in_img_array[25][9][9] <= img[11727];\
        in_img_array[25][9][10] <= img[11728];\
        in_img_array[25][9][11] <= img[11729];\
        in_img_array[25][9][12] <= img[11730];\
        in_img_array[25][9][13] <= img[11731];\
        in_img_array[25][9][14] <= img[11732];\
        in_img_array[25][9][15] <= img[11733];\
        in_img_array[25][9][16] <= img[11734];\
        in_img_array[25][9][17] <= img[11735];\
        in_img_array[25][10][0] <= img[11736];\
        in_img_array[25][10][1] <= img[11737];\
        in_img_array[25][10][2] <= img[11738];\
        in_img_array[25][10][3] <= img[11739];\
        in_img_array[25][10][4] <= img[11740];\
        in_img_array[25][10][5] <= img[11741];\
        in_img_array[25][10][6] <= img[11742];\
        in_img_array[25][10][7] <= img[11743];\
        in_img_array[25][10][8] <= img[11744];\
        in_img_array[25][10][9] <= img[11745];\
        in_img_array[25][10][10] <= img[11746];\
        in_img_array[25][10][11] <= img[11747];\
        in_img_array[25][10][12] <= img[11748];\
        in_img_array[25][10][13] <= img[11749];\
        in_img_array[25][10][14] <= img[11750];\
        in_img_array[25][10][15] <= img[11751];\
        in_img_array[25][10][16] <= img[11752];\
        in_img_array[25][10][17] <= img[11753];\
        in_img_array[25][11][0] <= img[11754];\
        in_img_array[25][11][1] <= img[11755];\
        in_img_array[25][11][2] <= img[11756];\
        in_img_array[25][11][3] <= img[11757];\
        in_img_array[25][11][4] <= img[11758];\
        in_img_array[25][11][5] <= img[11759];\
        in_img_array[25][11][6] <= img[11760];\
        in_img_array[25][11][7] <= img[11761];\
        in_img_array[25][11][8] <= img[11762];\
        in_img_array[25][11][9] <= img[11763];\
        in_img_array[25][11][10] <= img[11764];\
        in_img_array[25][11][11] <= img[11765];\
        in_img_array[25][11][12] <= img[11766];\
        in_img_array[25][11][13] <= img[11767];\
        in_img_array[25][11][14] <= img[11768];\
        in_img_array[25][11][15] <= img[11769];\
        in_img_array[25][11][16] <= img[11770];\
        in_img_array[25][11][17] <= img[11771];\
        in_img_array[25][12][0] <= img[11772];\
        in_img_array[25][12][1] <= img[11773];\
        in_img_array[25][12][2] <= img[11774];\
        in_img_array[25][12][3] <= img[11775];\
        in_img_array[25][12][4] <= img[11776];\
        in_img_array[25][12][5] <= img[11777];\
        in_img_array[25][12][6] <= img[11778];\
        in_img_array[25][12][7] <= img[11779];\
        in_img_array[25][12][8] <= img[11780];\
        in_img_array[25][12][9] <= img[11781];\
        in_img_array[25][12][10] <= img[11782];\
        in_img_array[25][12][11] <= img[11783];\
        in_img_array[25][12][12] <= img[11784];\
        in_img_array[25][12][13] <= img[11785];\
        in_img_array[25][12][14] <= img[11786];\
        in_img_array[25][12][15] <= img[11787];\
        in_img_array[25][12][16] <= img[11788];\
        in_img_array[25][12][17] <= img[11789];\
        in_img_array[25][13][0] <= img[11790];\
        in_img_array[25][13][1] <= img[11791];\
        in_img_array[25][13][2] <= img[11792];\
        in_img_array[25][13][3] <= img[11793];\
        in_img_array[25][13][4] <= img[11794];\
        in_img_array[25][13][5] <= img[11795];\
        in_img_array[25][13][6] <= img[11796];\
        in_img_array[25][13][7] <= img[11797];\
        in_img_array[25][13][8] <= img[11798];\
        in_img_array[25][13][9] <= img[11799];\
        in_img_array[25][13][10] <= img[11800];\
        in_img_array[25][13][11] <= img[11801];\
        in_img_array[25][13][12] <= img[11802];\
        in_img_array[25][13][13] <= img[11803];\
        in_img_array[25][13][14] <= img[11804];\
        in_img_array[25][13][15] <= img[11805];\
        in_img_array[25][13][16] <= img[11806];\
        in_img_array[25][13][17] <= img[11807];\
        in_img_array[25][14][0] <= img[11808];\
        in_img_array[25][14][1] <= img[11809];\
        in_img_array[25][14][2] <= img[11810];\
        in_img_array[25][14][3] <= img[11811];\
        in_img_array[25][14][4] <= img[11812];\
        in_img_array[25][14][5] <= img[11813];\
        in_img_array[25][14][6] <= img[11814];\
        in_img_array[25][14][7] <= img[11815];\
        in_img_array[25][14][8] <= img[11816];\
        in_img_array[25][14][9] <= img[11817];\
        in_img_array[25][14][10] <= img[11818];\
        in_img_array[25][14][11] <= img[11819];\
        in_img_array[25][14][12] <= img[11820];\
        in_img_array[25][14][13] <= img[11821];\
        in_img_array[25][14][14] <= img[11822];\
        in_img_array[25][14][15] <= img[11823];\
        in_img_array[25][14][16] <= img[11824];\
        in_img_array[25][14][17] <= img[11825];\
        in_img_array[25][15][0] <= img[11826];\
        in_img_array[25][15][1] <= img[11827];\
        in_img_array[25][15][2] <= img[11828];\
        in_img_array[25][15][3] <= img[11829];\
        in_img_array[25][15][4] <= img[11830];\
        in_img_array[25][15][5] <= img[11831];\
        in_img_array[25][15][6] <= img[11832];\
        in_img_array[25][15][7] <= img[11833];\
        in_img_array[25][15][8] <= img[11834];\
        in_img_array[25][15][9] <= img[11835];\
        in_img_array[25][15][10] <= img[11836];\
        in_img_array[25][15][11] <= img[11837];\
        in_img_array[25][15][12] <= img[11838];\
        in_img_array[25][15][13] <= img[11839];\
        in_img_array[25][15][14] <= img[11840];\
        in_img_array[25][15][15] <= img[11841];\
        in_img_array[25][15][16] <= img[11842];\
        in_img_array[25][15][17] <= img[11843];\
        in_img_array[25][16][0] <= img[11844];\
        in_img_array[25][16][1] <= img[11845];\
        in_img_array[25][16][2] <= img[11846];\
        in_img_array[25][16][3] <= img[11847];\
        in_img_array[25][16][4] <= img[11848];\
        in_img_array[25][16][5] <= img[11849];\
        in_img_array[25][16][6] <= img[11850];\
        in_img_array[25][16][7] <= img[11851];\
        in_img_array[25][16][8] <= img[11852];\
        in_img_array[25][16][9] <= img[11853];\
        in_img_array[25][16][10] <= img[11854];\
        in_img_array[25][16][11] <= img[11855];\
        in_img_array[25][16][12] <= img[11856];\
        in_img_array[25][16][13] <= img[11857];\
        in_img_array[25][16][14] <= img[11858];\
        in_img_array[25][16][15] <= img[11859];\
        in_img_array[25][16][16] <= img[11860];\
        in_img_array[25][16][17] <= img[11861];\
        in_img_array[25][17][0] <= img[11862];\
        in_img_array[25][17][1] <= img[11863];\
        in_img_array[25][17][2] <= img[11864];\
        in_img_array[25][17][3] <= img[11865];\
        in_img_array[25][17][4] <= img[11866];\
        in_img_array[25][17][5] <= img[11867];\
        in_img_array[25][17][6] <= img[11868];\
        in_img_array[25][17][7] <= img[11869];\
        in_img_array[25][17][8] <= img[11870];\
        in_img_array[25][17][9] <= img[11871];\
        in_img_array[25][17][10] <= img[11872];\
        in_img_array[25][17][11] <= img[11873];\
        in_img_array[25][17][12] <= img[11874];\
        in_img_array[25][17][13] <= img[11875];\
        in_img_array[25][17][14] <= img[11876];\
        in_img_array[25][17][15] <= img[11877];\
        in_img_array[25][17][16] <= img[11878];\
        in_img_array[25][17][17] <= img[11879];\
        in_img_array[25][18][0] <= img[11880];\
        in_img_array[25][18][1] <= img[11881];\
        in_img_array[25][18][2] <= img[11882];\
        in_img_array[25][18][3] <= img[11883];\
        in_img_array[25][18][4] <= img[11884];\
        in_img_array[25][18][5] <= img[11885];\
        in_img_array[25][18][6] <= img[11886];\
        in_img_array[25][18][7] <= img[11887];\
        in_img_array[25][18][8] <= img[11888];\
        in_img_array[25][18][9] <= img[11889];\
        in_img_array[25][18][10] <= img[11890];\
        in_img_array[25][18][11] <= img[11891];\
        in_img_array[25][18][12] <= img[11892];\
        in_img_array[25][18][13] <= img[11893];\
        in_img_array[25][18][14] <= img[11894];\
        in_img_array[25][18][15] <= img[11895];\
        in_img_array[25][18][16] <= img[11896];\
        in_img_array[25][18][17] <= img[11897];\
        in_img_array[25][19][0] <= img[11898];\
        in_img_array[25][19][1] <= img[11899];\
        in_img_array[25][19][2] <= img[11900];\
        in_img_array[25][19][3] <= img[11901];\
        in_img_array[25][19][4] <= img[11902];\
        in_img_array[25][19][5] <= img[11903];\
        in_img_array[25][19][6] <= img[11904];\
        in_img_array[25][19][7] <= img[11905];\
        in_img_array[25][19][8] <= img[11906];\
        in_img_array[25][19][9] <= img[11907];\
        in_img_array[25][19][10] <= img[11908];\
        in_img_array[25][19][11] <= img[11909];\
        in_img_array[25][19][12] <= img[11910];\
        in_img_array[25][19][13] <= img[11911];\
        in_img_array[25][19][14] <= img[11912];\
        in_img_array[25][19][15] <= img[11913];\
        in_img_array[25][19][16] <= img[11914];\
        in_img_array[25][19][17] <= img[11915];\
        in_img_array[25][20][0] <= img[11916];\
        in_img_array[25][20][1] <= img[11917];\
        in_img_array[25][20][2] <= img[11918];\
        in_img_array[25][20][3] <= img[11919];\
        in_img_array[25][20][4] <= img[11920];\
        in_img_array[25][20][5] <= img[11921];\
        in_img_array[25][20][6] <= img[11922];\
        in_img_array[25][20][7] <= img[11923];\
        in_img_array[25][20][8] <= img[11924];\
        in_img_array[25][20][9] <= img[11925];\
        in_img_array[25][20][10] <= img[11926];\
        in_img_array[25][20][11] <= img[11927];\
        in_img_array[25][20][12] <= img[11928];\
        in_img_array[25][20][13] <= img[11929];\
        in_img_array[25][20][14] <= img[11930];\
        in_img_array[25][20][15] <= img[11931];\
        in_img_array[25][20][16] <= img[11932];\
        in_img_array[25][20][17] <= img[11933];\
        in_img_array[25][21][0] <= img[11934];\
        in_img_array[25][21][1] <= img[11935];\
        in_img_array[25][21][2] <= img[11936];\
        in_img_array[25][21][3] <= img[11937];\
        in_img_array[25][21][4] <= img[11938];\
        in_img_array[25][21][5] <= img[11939];\
        in_img_array[25][21][6] <= img[11940];\
        in_img_array[25][21][7] <= img[11941];\
        in_img_array[25][21][8] <= img[11942];\
        in_img_array[25][21][9] <= img[11943];\
        in_img_array[25][21][10] <= img[11944];\
        in_img_array[25][21][11] <= img[11945];\
        in_img_array[25][21][12] <= img[11946];\
        in_img_array[25][21][13] <= img[11947];\
        in_img_array[25][21][14] <= img[11948];\
        in_img_array[25][21][15] <= img[11949];\
        in_img_array[25][21][16] <= img[11950];\
        in_img_array[25][21][17] <= img[11951];\
        in_img_array[25][22][0] <= img[11952];\
        in_img_array[25][22][1] <= img[11953];\
        in_img_array[25][22][2] <= img[11954];\
        in_img_array[25][22][3] <= img[11955];\
        in_img_array[25][22][4] <= img[11956];\
        in_img_array[25][22][5] <= img[11957];\
        in_img_array[25][22][6] <= img[11958];\
        in_img_array[25][22][7] <= img[11959];\
        in_img_array[25][22][8] <= img[11960];\
        in_img_array[25][22][9] <= img[11961];\
        in_img_array[25][22][10] <= img[11962];\
        in_img_array[25][22][11] <= img[11963];\
        in_img_array[25][22][12] <= img[11964];\
        in_img_array[25][22][13] <= img[11965];\
        in_img_array[25][22][14] <= img[11966];\
        in_img_array[25][22][15] <= img[11967];\
        in_img_array[25][22][16] <= img[11968];\
        in_img_array[25][22][17] <= img[11969];\
        in_img_array[25][23][0] <= img[11970];\
        in_img_array[25][23][1] <= img[11971];\
        in_img_array[25][23][2] <= img[11972];\
        in_img_array[25][23][3] <= img[11973];\
        in_img_array[25][23][4] <= img[11974];\
        in_img_array[25][23][5] <= img[11975];\
        in_img_array[25][23][6] <= img[11976];\
        in_img_array[25][23][7] <= img[11977];\
        in_img_array[25][23][8] <= img[11978];\
        in_img_array[25][23][9] <= img[11979];\
        in_img_array[25][23][10] <= img[11980];\
        in_img_array[25][23][11] <= img[11981];\
        in_img_array[25][23][12] <= img[11982];\
        in_img_array[25][23][13] <= img[11983];\
        in_img_array[25][23][14] <= img[11984];\
        in_img_array[25][23][15] <= img[11985];\
        in_img_array[25][23][16] <= img[11986];\
        in_img_array[25][23][17] <= img[11987];\
        in_img_array[25][24][0] <= img[11988];\
        in_img_array[25][24][1] <= img[11989];\
        in_img_array[25][24][2] <= img[11990];\
        in_img_array[25][24][3] <= img[11991];\
        in_img_array[25][24][4] <= img[11992];\
        in_img_array[25][24][5] <= img[11993];\
        in_img_array[25][24][6] <= img[11994];\
        in_img_array[25][24][7] <= img[11995];\
        in_img_array[25][24][8] <= img[11996];\
        in_img_array[25][24][9] <= img[11997];\
        in_img_array[25][24][10] <= img[11998];\
        in_img_array[25][24][11] <= img[11999];\
        in_img_array[25][24][12] <= img[12000];\
        in_img_array[25][24][13] <= img[12001];\
        in_img_array[25][24][14] <= img[12002];\
        in_img_array[25][24][15] <= img[12003];\
        in_img_array[25][24][16] <= img[12004];\
        in_img_array[25][24][17] <= img[12005];\
        in_img_array[25][25][0] <= img[12006];\
        in_img_array[25][25][1] <= img[12007];\
        in_img_array[25][25][2] <= img[12008];\
        in_img_array[25][25][3] <= img[12009];\
        in_img_array[25][25][4] <= img[12010];\
        in_img_array[25][25][5] <= img[12011];\
        in_img_array[25][25][6] <= img[12012];\
        in_img_array[25][25][7] <= img[12013];\
        in_img_array[25][25][8] <= img[12014];\
        in_img_array[25][25][9] <= img[12015];\
        in_img_array[25][25][10] <= img[12016];\
        in_img_array[25][25][11] <= img[12017];\
        in_img_array[25][25][12] <= img[12018];\
        in_img_array[25][25][13] <= img[12019];\
        in_img_array[25][25][14] <= img[12020];\
        in_img_array[25][25][15] <= img[12021];\
        in_img_array[25][25][16] <= img[12022];\
        in_img_array[25][25][17] <= img[12023];\
        in_img_array[25][26][0] <= img[12024];\
        in_img_array[25][26][1] <= img[12025];\
        in_img_array[25][26][2] <= img[12026];\
        in_img_array[25][26][3] <= img[12027];\
        in_img_array[25][26][4] <= img[12028];\
        in_img_array[25][26][5] <= img[12029];\
        in_img_array[25][26][6] <= img[12030];\
        in_img_array[25][26][7] <= img[12031];\
        in_img_array[25][26][8] <= img[12032];\
        in_img_array[25][26][9] <= img[12033];\
        in_img_array[25][26][10] <= img[12034];\
        in_img_array[25][26][11] <= img[12035];\
        in_img_array[25][26][12] <= img[12036];\
        in_img_array[25][26][13] <= img[12037];\
        in_img_array[25][26][14] <= img[12038];\
        in_img_array[25][26][15] <= img[12039];\
        in_img_array[25][26][16] <= img[12040];\
        in_img_array[25][26][17] <= img[12041];\
        in_img_array[25][27][0] <= img[12042];\
        in_img_array[25][27][1] <= img[12043];\
        in_img_array[25][27][2] <= img[12044];\
        in_img_array[25][27][3] <= img[12045];\
        in_img_array[25][27][4] <= img[12046];\
        in_img_array[25][27][5] <= img[12047];\
        in_img_array[25][27][6] <= img[12048];\
        in_img_array[25][27][7] <= img[12049];\
        in_img_array[25][27][8] <= img[12050];\
        in_img_array[25][27][9] <= img[12051];\
        in_img_array[25][27][10] <= img[12052];\
        in_img_array[25][27][11] <= img[12053];\
        in_img_array[25][27][12] <= img[12054];\
        in_img_array[25][27][13] <= img[12055];\
        in_img_array[25][27][14] <= img[12056];\
        in_img_array[25][27][15] <= img[12057];\
        in_img_array[25][27][16] <= img[12058];\
        in_img_array[25][27][17] <= img[12059];\
        in_img_array[25][28][0] <= img[12060];\
        in_img_array[25][28][1] <= img[12061];\
        in_img_array[25][28][2] <= img[12062];\
        in_img_array[25][28][3] <= img[12063];\
        in_img_array[25][28][4] <= img[12064];\
        in_img_array[25][28][5] <= img[12065];\
        in_img_array[25][28][6] <= img[12066];\
        in_img_array[25][28][7] <= img[12067];\
        in_img_array[25][28][8] <= img[12068];\
        in_img_array[25][28][9] <= img[12069];\
        in_img_array[25][28][10] <= img[12070];\
        in_img_array[25][28][11] <= img[12071];\
        in_img_array[25][28][12] <= img[12072];\
        in_img_array[25][28][13] <= img[12073];\
        in_img_array[25][28][14] <= img[12074];\
        in_img_array[25][28][15] <= img[12075];\
        in_img_array[25][28][16] <= img[12076];\
        in_img_array[25][28][17] <= img[12077];\
        in_img_array[25][29][0] <= img[12078];\
        in_img_array[25][29][1] <= img[12079];\
        in_img_array[25][29][2] <= img[12080];\
        in_img_array[25][29][3] <= img[12081];\
        in_img_array[25][29][4] <= img[12082];\
        in_img_array[25][29][5] <= img[12083];\
        in_img_array[25][29][6] <= img[12084];\
        in_img_array[25][29][7] <= img[12085];\
        in_img_array[25][29][8] <= img[12086];\
        in_img_array[25][29][9] <= img[12087];\
        in_img_array[25][29][10] <= img[12088];\
        in_img_array[25][29][11] <= img[12089];\
        in_img_array[25][29][12] <= img[12090];\
        in_img_array[25][29][13] <= img[12091];\
        in_img_array[25][29][14] <= img[12092];\
        in_img_array[25][29][15] <= img[12093];\
        in_img_array[25][29][16] <= img[12094];\
        in_img_array[25][29][17] <= img[12095];\
        in_img_array[26][2][0] <= img[12096];\
        in_img_array[26][2][1] <= img[12097];\
        in_img_array[26][2][2] <= img[12098];\
        in_img_array[26][2][3] <= img[12099];\
        in_img_array[26][2][4] <= img[12100];\
        in_img_array[26][2][5] <= img[12101];\
        in_img_array[26][2][6] <= img[12102];\
        in_img_array[26][2][7] <= img[12103];\
        in_img_array[26][2][8] <= img[12104];\
        in_img_array[26][2][9] <= img[12105];\
        in_img_array[26][2][10] <= img[12106];\
        in_img_array[26][2][11] <= img[12107];\
        in_img_array[26][2][12] <= img[12108];\
        in_img_array[26][2][13] <= img[12109];\
        in_img_array[26][2][14] <= img[12110];\
        in_img_array[26][2][15] <= img[12111];\
        in_img_array[26][2][16] <= img[12112];\
        in_img_array[26][2][17] <= img[12113];\
        in_img_array[26][3][0] <= img[12114];\
        in_img_array[26][3][1] <= img[12115];\
        in_img_array[26][3][2] <= img[12116];\
        in_img_array[26][3][3] <= img[12117];\
        in_img_array[26][3][4] <= img[12118];\
        in_img_array[26][3][5] <= img[12119];\
        in_img_array[26][3][6] <= img[12120];\
        in_img_array[26][3][7] <= img[12121];\
        in_img_array[26][3][8] <= img[12122];\
        in_img_array[26][3][9] <= img[12123];\
        in_img_array[26][3][10] <= img[12124];\
        in_img_array[26][3][11] <= img[12125];\
        in_img_array[26][3][12] <= img[12126];\
        in_img_array[26][3][13] <= img[12127];\
        in_img_array[26][3][14] <= img[12128];\
        in_img_array[26][3][15] <= img[12129];\
        in_img_array[26][3][16] <= img[12130];\
        in_img_array[26][3][17] <= img[12131];\
        in_img_array[26][4][0] <= img[12132];\
        in_img_array[26][4][1] <= img[12133];\
        in_img_array[26][4][2] <= img[12134];\
        in_img_array[26][4][3] <= img[12135];\
        in_img_array[26][4][4] <= img[12136];\
        in_img_array[26][4][5] <= img[12137];\
        in_img_array[26][4][6] <= img[12138];\
        in_img_array[26][4][7] <= img[12139];\
        in_img_array[26][4][8] <= img[12140];\
        in_img_array[26][4][9] <= img[12141];\
        in_img_array[26][4][10] <= img[12142];\
        in_img_array[26][4][11] <= img[12143];\
        in_img_array[26][4][12] <= img[12144];\
        in_img_array[26][4][13] <= img[12145];\
        in_img_array[26][4][14] <= img[12146];\
        in_img_array[26][4][15] <= img[12147];\
        in_img_array[26][4][16] <= img[12148];\
        in_img_array[26][4][17] <= img[12149];\
        in_img_array[26][5][0] <= img[12150];\
        in_img_array[26][5][1] <= img[12151];\
        in_img_array[26][5][2] <= img[12152];\
        in_img_array[26][5][3] <= img[12153];\
        in_img_array[26][5][4] <= img[12154];\
        in_img_array[26][5][5] <= img[12155];\
        in_img_array[26][5][6] <= img[12156];\
        in_img_array[26][5][7] <= img[12157];\
        in_img_array[26][5][8] <= img[12158];\
        in_img_array[26][5][9] <= img[12159];\
        in_img_array[26][5][10] <= img[12160];\
        in_img_array[26][5][11] <= img[12161];\
        in_img_array[26][5][12] <= img[12162];\
        in_img_array[26][5][13] <= img[12163];\
        in_img_array[26][5][14] <= img[12164];\
        in_img_array[26][5][15] <= img[12165];\
        in_img_array[26][5][16] <= img[12166];\
        in_img_array[26][5][17] <= img[12167];\
        in_img_array[26][6][0] <= img[12168];\
        in_img_array[26][6][1] <= img[12169];\
        in_img_array[26][6][2] <= img[12170];\
        in_img_array[26][6][3] <= img[12171];\
        in_img_array[26][6][4] <= img[12172];\
        in_img_array[26][6][5] <= img[12173];\
        in_img_array[26][6][6] <= img[12174];\
        in_img_array[26][6][7] <= img[12175];\
        in_img_array[26][6][8] <= img[12176];\
        in_img_array[26][6][9] <= img[12177];\
        in_img_array[26][6][10] <= img[12178];\
        in_img_array[26][6][11] <= img[12179];\
        in_img_array[26][6][12] <= img[12180];\
        in_img_array[26][6][13] <= img[12181];\
        in_img_array[26][6][14] <= img[12182];\
        in_img_array[26][6][15] <= img[12183];\
        in_img_array[26][6][16] <= img[12184];\
        in_img_array[26][6][17] <= img[12185];\
        in_img_array[26][7][0] <= img[12186];\
        in_img_array[26][7][1] <= img[12187];\
        in_img_array[26][7][2] <= img[12188];\
        in_img_array[26][7][3] <= img[12189];\
        in_img_array[26][7][4] <= img[12190];\
        in_img_array[26][7][5] <= img[12191];\
        in_img_array[26][7][6] <= img[12192];\
        in_img_array[26][7][7] <= img[12193];\
        in_img_array[26][7][8] <= img[12194];\
        in_img_array[26][7][9] <= img[12195];\
        in_img_array[26][7][10] <= img[12196];\
        in_img_array[26][7][11] <= img[12197];\
        in_img_array[26][7][12] <= img[12198];\
        in_img_array[26][7][13] <= img[12199];\
        in_img_array[26][7][14] <= img[12200];\
        in_img_array[26][7][15] <= img[12201];\
        in_img_array[26][7][16] <= img[12202];\
        in_img_array[26][7][17] <= img[12203];\
        in_img_array[26][8][0] <= img[12204];\
        in_img_array[26][8][1] <= img[12205];\
        in_img_array[26][8][2] <= img[12206];\
        in_img_array[26][8][3] <= img[12207];\
        in_img_array[26][8][4] <= img[12208];\
        in_img_array[26][8][5] <= img[12209];\
        in_img_array[26][8][6] <= img[12210];\
        in_img_array[26][8][7] <= img[12211];\
        in_img_array[26][8][8] <= img[12212];\
        in_img_array[26][8][9] <= img[12213];\
        in_img_array[26][8][10] <= img[12214];\
        in_img_array[26][8][11] <= img[12215];\
        in_img_array[26][8][12] <= img[12216];\
        in_img_array[26][8][13] <= img[12217];\
        in_img_array[26][8][14] <= img[12218];\
        in_img_array[26][8][15] <= img[12219];\
        in_img_array[26][8][16] <= img[12220];\
        in_img_array[26][8][17] <= img[12221];\
        in_img_array[26][9][0] <= img[12222];\
        in_img_array[26][9][1] <= img[12223];\
        in_img_array[26][9][2] <= img[12224];\
        in_img_array[26][9][3] <= img[12225];\
        in_img_array[26][9][4] <= img[12226];\
        in_img_array[26][9][5] <= img[12227];\
        in_img_array[26][9][6] <= img[12228];\
        in_img_array[26][9][7] <= img[12229];\
        in_img_array[26][9][8] <= img[12230];\
        in_img_array[26][9][9] <= img[12231];\
        in_img_array[26][9][10] <= img[12232];\
        in_img_array[26][9][11] <= img[12233];\
        in_img_array[26][9][12] <= img[12234];\
        in_img_array[26][9][13] <= img[12235];\
        in_img_array[26][9][14] <= img[12236];\
        in_img_array[26][9][15] <= img[12237];\
        in_img_array[26][9][16] <= img[12238];\
        in_img_array[26][9][17] <= img[12239];\
        in_img_array[26][10][0] <= img[12240];\
        in_img_array[26][10][1] <= img[12241];\
        in_img_array[26][10][2] <= img[12242];\
        in_img_array[26][10][3] <= img[12243];\
        in_img_array[26][10][4] <= img[12244];\
        in_img_array[26][10][5] <= img[12245];\
        in_img_array[26][10][6] <= img[12246];\
        in_img_array[26][10][7] <= img[12247];\
        in_img_array[26][10][8] <= img[12248];\
        in_img_array[26][10][9] <= img[12249];\
        in_img_array[26][10][10] <= img[12250];\
        in_img_array[26][10][11] <= img[12251];\
        in_img_array[26][10][12] <= img[12252];\
        in_img_array[26][10][13] <= img[12253];\
        in_img_array[26][10][14] <= img[12254];\
        in_img_array[26][10][15] <= img[12255];\
        in_img_array[26][10][16] <= img[12256];\
        in_img_array[26][10][17] <= img[12257];\
        in_img_array[26][11][0] <= img[12258];\
        in_img_array[26][11][1] <= img[12259];\
        in_img_array[26][11][2] <= img[12260];\
        in_img_array[26][11][3] <= img[12261];\
        in_img_array[26][11][4] <= img[12262];\
        in_img_array[26][11][5] <= img[12263];\
        in_img_array[26][11][6] <= img[12264];\
        in_img_array[26][11][7] <= img[12265];\
        in_img_array[26][11][8] <= img[12266];\
        in_img_array[26][11][9] <= img[12267];\
        in_img_array[26][11][10] <= img[12268];\
        in_img_array[26][11][11] <= img[12269];\
        in_img_array[26][11][12] <= img[12270];\
        in_img_array[26][11][13] <= img[12271];\
        in_img_array[26][11][14] <= img[12272];\
        in_img_array[26][11][15] <= img[12273];\
        in_img_array[26][11][16] <= img[12274];\
        in_img_array[26][11][17] <= img[12275];\
        in_img_array[26][12][0] <= img[12276];\
        in_img_array[26][12][1] <= img[12277];\
        in_img_array[26][12][2] <= img[12278];\
        in_img_array[26][12][3] <= img[12279];\
        in_img_array[26][12][4] <= img[12280];\
        in_img_array[26][12][5] <= img[12281];\
        in_img_array[26][12][6] <= img[12282];\
        in_img_array[26][12][7] <= img[12283];\
        in_img_array[26][12][8] <= img[12284];\
        in_img_array[26][12][9] <= img[12285];\
        in_img_array[26][12][10] <= img[12286];\
        in_img_array[26][12][11] <= img[12287];\
        in_img_array[26][12][12] <= img[12288];\
        in_img_array[26][12][13] <= img[12289];\
        in_img_array[26][12][14] <= img[12290];\
        in_img_array[26][12][15] <= img[12291];\
        in_img_array[26][12][16] <= img[12292];\
        in_img_array[26][12][17] <= img[12293];\
        in_img_array[26][13][0] <= img[12294];\
        in_img_array[26][13][1] <= img[12295];\
        in_img_array[26][13][2] <= img[12296];\
        in_img_array[26][13][3] <= img[12297];\
        in_img_array[26][13][4] <= img[12298];\
        in_img_array[26][13][5] <= img[12299];\
        in_img_array[26][13][6] <= img[12300];\
        in_img_array[26][13][7] <= img[12301];\
        in_img_array[26][13][8] <= img[12302];\
        in_img_array[26][13][9] <= img[12303];\
        in_img_array[26][13][10] <= img[12304];\
        in_img_array[26][13][11] <= img[12305];\
        in_img_array[26][13][12] <= img[12306];\
        in_img_array[26][13][13] <= img[12307];\
        in_img_array[26][13][14] <= img[12308];\
        in_img_array[26][13][15] <= img[12309];\
        in_img_array[26][13][16] <= img[12310];\
        in_img_array[26][13][17] <= img[12311];\
        in_img_array[26][14][0] <= img[12312];\
        in_img_array[26][14][1] <= img[12313];\
        in_img_array[26][14][2] <= img[12314];\
        in_img_array[26][14][3] <= img[12315];\
        in_img_array[26][14][4] <= img[12316];\
        in_img_array[26][14][5] <= img[12317];\
        in_img_array[26][14][6] <= img[12318];\
        in_img_array[26][14][7] <= img[12319];\
        in_img_array[26][14][8] <= img[12320];\
        in_img_array[26][14][9] <= img[12321];\
        in_img_array[26][14][10] <= img[12322];\
        in_img_array[26][14][11] <= img[12323];\
        in_img_array[26][14][12] <= img[12324];\
        in_img_array[26][14][13] <= img[12325];\
        in_img_array[26][14][14] <= img[12326];\
        in_img_array[26][14][15] <= img[12327];\
        in_img_array[26][14][16] <= img[12328];\
        in_img_array[26][14][17] <= img[12329];\
        in_img_array[26][15][0] <= img[12330];\
        in_img_array[26][15][1] <= img[12331];\
        in_img_array[26][15][2] <= img[12332];\
        in_img_array[26][15][3] <= img[12333];\
        in_img_array[26][15][4] <= img[12334];\
        in_img_array[26][15][5] <= img[12335];\
        in_img_array[26][15][6] <= img[12336];\
        in_img_array[26][15][7] <= img[12337];\
        in_img_array[26][15][8] <= img[12338];\
        in_img_array[26][15][9] <= img[12339];\
        in_img_array[26][15][10] <= img[12340];\
        in_img_array[26][15][11] <= img[12341];\
        in_img_array[26][15][12] <= img[12342];\
        in_img_array[26][15][13] <= img[12343];\
        in_img_array[26][15][14] <= img[12344];\
        in_img_array[26][15][15] <= img[12345];\
        in_img_array[26][15][16] <= img[12346];\
        in_img_array[26][15][17] <= img[12347];\
        in_img_array[26][16][0] <= img[12348];\
        in_img_array[26][16][1] <= img[12349];\
        in_img_array[26][16][2] <= img[12350];\
        in_img_array[26][16][3] <= img[12351];\
        in_img_array[26][16][4] <= img[12352];\
        in_img_array[26][16][5] <= img[12353];\
        in_img_array[26][16][6] <= img[12354];\
        in_img_array[26][16][7] <= img[12355];\
        in_img_array[26][16][8] <= img[12356];\
        in_img_array[26][16][9] <= img[12357];\
        in_img_array[26][16][10] <= img[12358];\
        in_img_array[26][16][11] <= img[12359];\
        in_img_array[26][16][12] <= img[12360];\
        in_img_array[26][16][13] <= img[12361];\
        in_img_array[26][16][14] <= img[12362];\
        in_img_array[26][16][15] <= img[12363];\
        in_img_array[26][16][16] <= img[12364];\
        in_img_array[26][16][17] <= img[12365];\
        in_img_array[26][17][0] <= img[12366];\
        in_img_array[26][17][1] <= img[12367];\
        in_img_array[26][17][2] <= img[12368];\
        in_img_array[26][17][3] <= img[12369];\
        in_img_array[26][17][4] <= img[12370];\
        in_img_array[26][17][5] <= img[12371];\
        in_img_array[26][17][6] <= img[12372];\
        in_img_array[26][17][7] <= img[12373];\
        in_img_array[26][17][8] <= img[12374];\
        in_img_array[26][17][9] <= img[12375];\
        in_img_array[26][17][10] <= img[12376];\
        in_img_array[26][17][11] <= img[12377];\
        in_img_array[26][17][12] <= img[12378];\
        in_img_array[26][17][13] <= img[12379];\
        in_img_array[26][17][14] <= img[12380];\
        in_img_array[26][17][15] <= img[12381];\
        in_img_array[26][17][16] <= img[12382];\
        in_img_array[26][17][17] <= img[12383];\
        in_img_array[26][18][0] <= img[12384];\
        in_img_array[26][18][1] <= img[12385];\
        in_img_array[26][18][2] <= img[12386];\
        in_img_array[26][18][3] <= img[12387];\
        in_img_array[26][18][4] <= img[12388];\
        in_img_array[26][18][5] <= img[12389];\
        in_img_array[26][18][6] <= img[12390];\
        in_img_array[26][18][7] <= img[12391];\
        in_img_array[26][18][8] <= img[12392];\
        in_img_array[26][18][9] <= img[12393];\
        in_img_array[26][18][10] <= img[12394];\
        in_img_array[26][18][11] <= img[12395];\
        in_img_array[26][18][12] <= img[12396];\
        in_img_array[26][18][13] <= img[12397];\
        in_img_array[26][18][14] <= img[12398];\
        in_img_array[26][18][15] <= img[12399];\
        in_img_array[26][18][16] <= img[12400];\
        in_img_array[26][18][17] <= img[12401];\
        in_img_array[26][19][0] <= img[12402];\
        in_img_array[26][19][1] <= img[12403];\
        in_img_array[26][19][2] <= img[12404];\
        in_img_array[26][19][3] <= img[12405];\
        in_img_array[26][19][4] <= img[12406];\
        in_img_array[26][19][5] <= img[12407];\
        in_img_array[26][19][6] <= img[12408];\
        in_img_array[26][19][7] <= img[12409];\
        in_img_array[26][19][8] <= img[12410];\
        in_img_array[26][19][9] <= img[12411];\
        in_img_array[26][19][10] <= img[12412];\
        in_img_array[26][19][11] <= img[12413];\
        in_img_array[26][19][12] <= img[12414];\
        in_img_array[26][19][13] <= img[12415];\
        in_img_array[26][19][14] <= img[12416];\
        in_img_array[26][19][15] <= img[12417];\
        in_img_array[26][19][16] <= img[12418];\
        in_img_array[26][19][17] <= img[12419];\
        in_img_array[26][20][0] <= img[12420];\
        in_img_array[26][20][1] <= img[12421];\
        in_img_array[26][20][2] <= img[12422];\
        in_img_array[26][20][3] <= img[12423];\
        in_img_array[26][20][4] <= img[12424];\
        in_img_array[26][20][5] <= img[12425];\
        in_img_array[26][20][6] <= img[12426];\
        in_img_array[26][20][7] <= img[12427];\
        in_img_array[26][20][8] <= img[12428];\
        in_img_array[26][20][9] <= img[12429];\
        in_img_array[26][20][10] <= img[12430];\
        in_img_array[26][20][11] <= img[12431];\
        in_img_array[26][20][12] <= img[12432];\
        in_img_array[26][20][13] <= img[12433];\
        in_img_array[26][20][14] <= img[12434];\
        in_img_array[26][20][15] <= img[12435];\
        in_img_array[26][20][16] <= img[12436];\
        in_img_array[26][20][17] <= img[12437];\
        in_img_array[26][21][0] <= img[12438];\
        in_img_array[26][21][1] <= img[12439];\
        in_img_array[26][21][2] <= img[12440];\
        in_img_array[26][21][3] <= img[12441];\
        in_img_array[26][21][4] <= img[12442];\
        in_img_array[26][21][5] <= img[12443];\
        in_img_array[26][21][6] <= img[12444];\
        in_img_array[26][21][7] <= img[12445];\
        in_img_array[26][21][8] <= img[12446];\
        in_img_array[26][21][9] <= img[12447];\
        in_img_array[26][21][10] <= img[12448];\
        in_img_array[26][21][11] <= img[12449];\
        in_img_array[26][21][12] <= img[12450];\
        in_img_array[26][21][13] <= img[12451];\
        in_img_array[26][21][14] <= img[12452];\
        in_img_array[26][21][15] <= img[12453];\
        in_img_array[26][21][16] <= img[12454];\
        in_img_array[26][21][17] <= img[12455];\
        in_img_array[26][22][0] <= img[12456];\
        in_img_array[26][22][1] <= img[12457];\
        in_img_array[26][22][2] <= img[12458];\
        in_img_array[26][22][3] <= img[12459];\
        in_img_array[26][22][4] <= img[12460];\
        in_img_array[26][22][5] <= img[12461];\
        in_img_array[26][22][6] <= img[12462];\
        in_img_array[26][22][7] <= img[12463];\
        in_img_array[26][22][8] <= img[12464];\
        in_img_array[26][22][9] <= img[12465];\
        in_img_array[26][22][10] <= img[12466];\
        in_img_array[26][22][11] <= img[12467];\
        in_img_array[26][22][12] <= img[12468];\
        in_img_array[26][22][13] <= img[12469];\
        in_img_array[26][22][14] <= img[12470];\
        in_img_array[26][22][15] <= img[12471];\
        in_img_array[26][22][16] <= img[12472];\
        in_img_array[26][22][17] <= img[12473];\
        in_img_array[26][23][0] <= img[12474];\
        in_img_array[26][23][1] <= img[12475];\
        in_img_array[26][23][2] <= img[12476];\
        in_img_array[26][23][3] <= img[12477];\
        in_img_array[26][23][4] <= img[12478];\
        in_img_array[26][23][5] <= img[12479];\
        in_img_array[26][23][6] <= img[12480];\
        in_img_array[26][23][7] <= img[12481];\
        in_img_array[26][23][8] <= img[12482];\
        in_img_array[26][23][9] <= img[12483];\
        in_img_array[26][23][10] <= img[12484];\
        in_img_array[26][23][11] <= img[12485];\
        in_img_array[26][23][12] <= img[12486];\
        in_img_array[26][23][13] <= img[12487];\
        in_img_array[26][23][14] <= img[12488];\
        in_img_array[26][23][15] <= img[12489];\
        in_img_array[26][23][16] <= img[12490];\
        in_img_array[26][23][17] <= img[12491];\
        in_img_array[26][24][0] <= img[12492];\
        in_img_array[26][24][1] <= img[12493];\
        in_img_array[26][24][2] <= img[12494];\
        in_img_array[26][24][3] <= img[12495];\
        in_img_array[26][24][4] <= img[12496];\
        in_img_array[26][24][5] <= img[12497];\
        in_img_array[26][24][6] <= img[12498];\
        in_img_array[26][24][7] <= img[12499];\
        in_img_array[26][24][8] <= img[12500];\
        in_img_array[26][24][9] <= img[12501];\
        in_img_array[26][24][10] <= img[12502];\
        in_img_array[26][24][11] <= img[12503];\
        in_img_array[26][24][12] <= img[12504];\
        in_img_array[26][24][13] <= img[12505];\
        in_img_array[26][24][14] <= img[12506];\
        in_img_array[26][24][15] <= img[12507];\
        in_img_array[26][24][16] <= img[12508];\
        in_img_array[26][24][17] <= img[12509];\
        in_img_array[26][25][0] <= img[12510];\
        in_img_array[26][25][1] <= img[12511];\
        in_img_array[26][25][2] <= img[12512];\
        in_img_array[26][25][3] <= img[12513];\
        in_img_array[26][25][4] <= img[12514];\
        in_img_array[26][25][5] <= img[12515];\
        in_img_array[26][25][6] <= img[12516];\
        in_img_array[26][25][7] <= img[12517];\
        in_img_array[26][25][8] <= img[12518];\
        in_img_array[26][25][9] <= img[12519];\
        in_img_array[26][25][10] <= img[12520];\
        in_img_array[26][25][11] <= img[12521];\
        in_img_array[26][25][12] <= img[12522];\
        in_img_array[26][25][13] <= img[12523];\
        in_img_array[26][25][14] <= img[12524];\
        in_img_array[26][25][15] <= img[12525];\
        in_img_array[26][25][16] <= img[12526];\
        in_img_array[26][25][17] <= img[12527];\
        in_img_array[26][26][0] <= img[12528];\
        in_img_array[26][26][1] <= img[12529];\
        in_img_array[26][26][2] <= img[12530];\
        in_img_array[26][26][3] <= img[12531];\
        in_img_array[26][26][4] <= img[12532];\
        in_img_array[26][26][5] <= img[12533];\
        in_img_array[26][26][6] <= img[12534];\
        in_img_array[26][26][7] <= img[12535];\
        in_img_array[26][26][8] <= img[12536];\
        in_img_array[26][26][9] <= img[12537];\
        in_img_array[26][26][10] <= img[12538];\
        in_img_array[26][26][11] <= img[12539];\
        in_img_array[26][26][12] <= img[12540];\
        in_img_array[26][26][13] <= img[12541];\
        in_img_array[26][26][14] <= img[12542];\
        in_img_array[26][26][15] <= img[12543];\
        in_img_array[26][26][16] <= img[12544];\
        in_img_array[26][26][17] <= img[12545];\
        in_img_array[26][27][0] <= img[12546];\
        in_img_array[26][27][1] <= img[12547];\
        in_img_array[26][27][2] <= img[12548];\
        in_img_array[26][27][3] <= img[12549];\
        in_img_array[26][27][4] <= img[12550];\
        in_img_array[26][27][5] <= img[12551];\
        in_img_array[26][27][6] <= img[12552];\
        in_img_array[26][27][7] <= img[12553];\
        in_img_array[26][27][8] <= img[12554];\
        in_img_array[26][27][9] <= img[12555];\
        in_img_array[26][27][10] <= img[12556];\
        in_img_array[26][27][11] <= img[12557];\
        in_img_array[26][27][12] <= img[12558];\
        in_img_array[26][27][13] <= img[12559];\
        in_img_array[26][27][14] <= img[12560];\
        in_img_array[26][27][15] <= img[12561];\
        in_img_array[26][27][16] <= img[12562];\
        in_img_array[26][27][17] <= img[12563];\
        in_img_array[26][28][0] <= img[12564];\
        in_img_array[26][28][1] <= img[12565];\
        in_img_array[26][28][2] <= img[12566];\
        in_img_array[26][28][3] <= img[12567];\
        in_img_array[26][28][4] <= img[12568];\
        in_img_array[26][28][5] <= img[12569];\
        in_img_array[26][28][6] <= img[12570];\
        in_img_array[26][28][7] <= img[12571];\
        in_img_array[26][28][8] <= img[12572];\
        in_img_array[26][28][9] <= img[12573];\
        in_img_array[26][28][10] <= img[12574];\
        in_img_array[26][28][11] <= img[12575];\
        in_img_array[26][28][12] <= img[12576];\
        in_img_array[26][28][13] <= img[12577];\
        in_img_array[26][28][14] <= img[12578];\
        in_img_array[26][28][15] <= img[12579];\
        in_img_array[26][28][16] <= img[12580];\
        in_img_array[26][28][17] <= img[12581];\
        in_img_array[26][29][0] <= img[12582];\
        in_img_array[26][29][1] <= img[12583];\
        in_img_array[26][29][2] <= img[12584];\
        in_img_array[26][29][3] <= img[12585];\
        in_img_array[26][29][4] <= img[12586];\
        in_img_array[26][29][5] <= img[12587];\
        in_img_array[26][29][6] <= img[12588];\
        in_img_array[26][29][7] <= img[12589];\
        in_img_array[26][29][8] <= img[12590];\
        in_img_array[26][29][9] <= img[12591];\
        in_img_array[26][29][10] <= img[12592];\
        in_img_array[26][29][11] <= img[12593];\
        in_img_array[26][29][12] <= img[12594];\
        in_img_array[26][29][13] <= img[12595];\
        in_img_array[26][29][14] <= img[12596];\
        in_img_array[26][29][15] <= img[12597];\
        in_img_array[26][29][16] <= img[12598];\
        in_img_array[26][29][17] <= img[12599];\
        in_img_array[27][2][0] <= img[12600];\
        in_img_array[27][2][1] <= img[12601];\
        in_img_array[27][2][2] <= img[12602];\
        in_img_array[27][2][3] <= img[12603];\
        in_img_array[27][2][4] <= img[12604];\
        in_img_array[27][2][5] <= img[12605];\
        in_img_array[27][2][6] <= img[12606];\
        in_img_array[27][2][7] <= img[12607];\
        in_img_array[27][2][8] <= img[12608];\
        in_img_array[27][2][9] <= img[12609];\
        in_img_array[27][2][10] <= img[12610];\
        in_img_array[27][2][11] <= img[12611];\
        in_img_array[27][2][12] <= img[12612];\
        in_img_array[27][2][13] <= img[12613];\
        in_img_array[27][2][14] <= img[12614];\
        in_img_array[27][2][15] <= img[12615];\
        in_img_array[27][2][16] <= img[12616];\
        in_img_array[27][2][17] <= img[12617];\
        in_img_array[27][3][0] <= img[12618];\
        in_img_array[27][3][1] <= img[12619];\
        in_img_array[27][3][2] <= img[12620];\
        in_img_array[27][3][3] <= img[12621];\
        in_img_array[27][3][4] <= img[12622];\
        in_img_array[27][3][5] <= img[12623];\
        in_img_array[27][3][6] <= img[12624];\
        in_img_array[27][3][7] <= img[12625];\
        in_img_array[27][3][8] <= img[12626];\
        in_img_array[27][3][9] <= img[12627];\
        in_img_array[27][3][10] <= img[12628];\
        in_img_array[27][3][11] <= img[12629];\
        in_img_array[27][3][12] <= img[12630];\
        in_img_array[27][3][13] <= img[12631];\
        in_img_array[27][3][14] <= img[12632];\
        in_img_array[27][3][15] <= img[12633];\
        in_img_array[27][3][16] <= img[12634];\
        in_img_array[27][3][17] <= img[12635];\
        in_img_array[27][4][0] <= img[12636];\
        in_img_array[27][4][1] <= img[12637];\
        in_img_array[27][4][2] <= img[12638];\
        in_img_array[27][4][3] <= img[12639];\
        in_img_array[27][4][4] <= img[12640];\
        in_img_array[27][4][5] <= img[12641];\
        in_img_array[27][4][6] <= img[12642];\
        in_img_array[27][4][7] <= img[12643];\
        in_img_array[27][4][8] <= img[12644];\
        in_img_array[27][4][9] <= img[12645];\
        in_img_array[27][4][10] <= img[12646];\
        in_img_array[27][4][11] <= img[12647];\
        in_img_array[27][4][12] <= img[12648];\
        in_img_array[27][4][13] <= img[12649];\
        in_img_array[27][4][14] <= img[12650];\
        in_img_array[27][4][15] <= img[12651];\
        in_img_array[27][4][16] <= img[12652];\
        in_img_array[27][4][17] <= img[12653];\
        in_img_array[27][5][0] <= img[12654];\
        in_img_array[27][5][1] <= img[12655];\
        in_img_array[27][5][2] <= img[12656];\
        in_img_array[27][5][3] <= img[12657];\
        in_img_array[27][5][4] <= img[12658];\
        in_img_array[27][5][5] <= img[12659];\
        in_img_array[27][5][6] <= img[12660];\
        in_img_array[27][5][7] <= img[12661];\
        in_img_array[27][5][8] <= img[12662];\
        in_img_array[27][5][9] <= img[12663];\
        in_img_array[27][5][10] <= img[12664];\
        in_img_array[27][5][11] <= img[12665];\
        in_img_array[27][5][12] <= img[12666];\
        in_img_array[27][5][13] <= img[12667];\
        in_img_array[27][5][14] <= img[12668];\
        in_img_array[27][5][15] <= img[12669];\
        in_img_array[27][5][16] <= img[12670];\
        in_img_array[27][5][17] <= img[12671];\
        in_img_array[27][6][0] <= img[12672];\
        in_img_array[27][6][1] <= img[12673];\
        in_img_array[27][6][2] <= img[12674];\
        in_img_array[27][6][3] <= img[12675];\
        in_img_array[27][6][4] <= img[12676];\
        in_img_array[27][6][5] <= img[12677];\
        in_img_array[27][6][6] <= img[12678];\
        in_img_array[27][6][7] <= img[12679];\
        in_img_array[27][6][8] <= img[12680];\
        in_img_array[27][6][9] <= img[12681];\
        in_img_array[27][6][10] <= img[12682];\
        in_img_array[27][6][11] <= img[12683];\
        in_img_array[27][6][12] <= img[12684];\
        in_img_array[27][6][13] <= img[12685];\
        in_img_array[27][6][14] <= img[12686];\
        in_img_array[27][6][15] <= img[12687];\
        in_img_array[27][6][16] <= img[12688];\
        in_img_array[27][6][17] <= img[12689];\
        in_img_array[27][7][0] <= img[12690];\
        in_img_array[27][7][1] <= img[12691];\
        in_img_array[27][7][2] <= img[12692];\
        in_img_array[27][7][3] <= img[12693];\
        in_img_array[27][7][4] <= img[12694];\
        in_img_array[27][7][5] <= img[12695];\
        in_img_array[27][7][6] <= img[12696];\
        in_img_array[27][7][7] <= img[12697];\
        in_img_array[27][7][8] <= img[12698];\
        in_img_array[27][7][9] <= img[12699];\
        in_img_array[27][7][10] <= img[12700];\
        in_img_array[27][7][11] <= img[12701];\
        in_img_array[27][7][12] <= img[12702];\
        in_img_array[27][7][13] <= img[12703];\
        in_img_array[27][7][14] <= img[12704];\
        in_img_array[27][7][15] <= img[12705];\
        in_img_array[27][7][16] <= img[12706];\
        in_img_array[27][7][17] <= img[12707];\
        in_img_array[27][8][0] <= img[12708];\
        in_img_array[27][8][1] <= img[12709];\
        in_img_array[27][8][2] <= img[12710];\
        in_img_array[27][8][3] <= img[12711];\
        in_img_array[27][8][4] <= img[12712];\
        in_img_array[27][8][5] <= img[12713];\
        in_img_array[27][8][6] <= img[12714];\
        in_img_array[27][8][7] <= img[12715];\
        in_img_array[27][8][8] <= img[12716];\
        in_img_array[27][8][9] <= img[12717];\
        in_img_array[27][8][10] <= img[12718];\
        in_img_array[27][8][11] <= img[12719];\
        in_img_array[27][8][12] <= img[12720];\
        in_img_array[27][8][13] <= img[12721];\
        in_img_array[27][8][14] <= img[12722];\
        in_img_array[27][8][15] <= img[12723];\
        in_img_array[27][8][16] <= img[12724];\
        in_img_array[27][8][17] <= img[12725];\
        in_img_array[27][9][0] <= img[12726];\
        in_img_array[27][9][1] <= img[12727];\
        in_img_array[27][9][2] <= img[12728];\
        in_img_array[27][9][3] <= img[12729];\
        in_img_array[27][9][4] <= img[12730];\
        in_img_array[27][9][5] <= img[12731];\
        in_img_array[27][9][6] <= img[12732];\
        in_img_array[27][9][7] <= img[12733];\
        in_img_array[27][9][8] <= img[12734];\
        in_img_array[27][9][9] <= img[12735];\
        in_img_array[27][9][10] <= img[12736];\
        in_img_array[27][9][11] <= img[12737];\
        in_img_array[27][9][12] <= img[12738];\
        in_img_array[27][9][13] <= img[12739];\
        in_img_array[27][9][14] <= img[12740];\
        in_img_array[27][9][15] <= img[12741];\
        in_img_array[27][9][16] <= img[12742];\
        in_img_array[27][9][17] <= img[12743];\
        in_img_array[27][10][0] <= img[12744];\
        in_img_array[27][10][1] <= img[12745];\
        in_img_array[27][10][2] <= img[12746];\
        in_img_array[27][10][3] <= img[12747];\
        in_img_array[27][10][4] <= img[12748];\
        in_img_array[27][10][5] <= img[12749];\
        in_img_array[27][10][6] <= img[12750];\
        in_img_array[27][10][7] <= img[12751];\
        in_img_array[27][10][8] <= img[12752];\
        in_img_array[27][10][9] <= img[12753];\
        in_img_array[27][10][10] <= img[12754];\
        in_img_array[27][10][11] <= img[12755];\
        in_img_array[27][10][12] <= img[12756];\
        in_img_array[27][10][13] <= img[12757];\
        in_img_array[27][10][14] <= img[12758];\
        in_img_array[27][10][15] <= img[12759];\
        in_img_array[27][10][16] <= img[12760];\
        in_img_array[27][10][17] <= img[12761];\
        in_img_array[27][11][0] <= img[12762];\
        in_img_array[27][11][1] <= img[12763];\
        in_img_array[27][11][2] <= img[12764];\
        in_img_array[27][11][3] <= img[12765];\
        in_img_array[27][11][4] <= img[12766];\
        in_img_array[27][11][5] <= img[12767];\
        in_img_array[27][11][6] <= img[12768];\
        in_img_array[27][11][7] <= img[12769];\
        in_img_array[27][11][8] <= img[12770];\
        in_img_array[27][11][9] <= img[12771];\
        in_img_array[27][11][10] <= img[12772];\
        in_img_array[27][11][11] <= img[12773];\
        in_img_array[27][11][12] <= img[12774];\
        in_img_array[27][11][13] <= img[12775];\
        in_img_array[27][11][14] <= img[12776];\
        in_img_array[27][11][15] <= img[12777];\
        in_img_array[27][11][16] <= img[12778];\
        in_img_array[27][11][17] <= img[12779];\
        in_img_array[27][12][0] <= img[12780];\
        in_img_array[27][12][1] <= img[12781];\
        in_img_array[27][12][2] <= img[12782];\
        in_img_array[27][12][3] <= img[12783];\
        in_img_array[27][12][4] <= img[12784];\
        in_img_array[27][12][5] <= img[12785];\
        in_img_array[27][12][6] <= img[12786];\
        in_img_array[27][12][7] <= img[12787];\
        in_img_array[27][12][8] <= img[12788];\
        in_img_array[27][12][9] <= img[12789];\
        in_img_array[27][12][10] <= img[12790];\
        in_img_array[27][12][11] <= img[12791];\
        in_img_array[27][12][12] <= img[12792];\
        in_img_array[27][12][13] <= img[12793];\
        in_img_array[27][12][14] <= img[12794];\
        in_img_array[27][12][15] <= img[12795];\
        in_img_array[27][12][16] <= img[12796];\
        in_img_array[27][12][17] <= img[12797];\
        in_img_array[27][13][0] <= img[12798];\
        in_img_array[27][13][1] <= img[12799];\
        in_img_array[27][13][2] <= img[12800];\
        in_img_array[27][13][3] <= img[12801];\
        in_img_array[27][13][4] <= img[12802];\
        in_img_array[27][13][5] <= img[12803];\
        in_img_array[27][13][6] <= img[12804];\
        in_img_array[27][13][7] <= img[12805];\
        in_img_array[27][13][8] <= img[12806];\
        in_img_array[27][13][9] <= img[12807];\
        in_img_array[27][13][10] <= img[12808];\
        in_img_array[27][13][11] <= img[12809];\
        in_img_array[27][13][12] <= img[12810];\
        in_img_array[27][13][13] <= img[12811];\
        in_img_array[27][13][14] <= img[12812];\
        in_img_array[27][13][15] <= img[12813];\
        in_img_array[27][13][16] <= img[12814];\
        in_img_array[27][13][17] <= img[12815];\
        in_img_array[27][14][0] <= img[12816];\
        in_img_array[27][14][1] <= img[12817];\
        in_img_array[27][14][2] <= img[12818];\
        in_img_array[27][14][3] <= img[12819];\
        in_img_array[27][14][4] <= img[12820];\
        in_img_array[27][14][5] <= img[12821];\
        in_img_array[27][14][6] <= img[12822];\
        in_img_array[27][14][7] <= img[12823];\
        in_img_array[27][14][8] <= img[12824];\
        in_img_array[27][14][9] <= img[12825];\
        in_img_array[27][14][10] <= img[12826];\
        in_img_array[27][14][11] <= img[12827];\
        in_img_array[27][14][12] <= img[12828];\
        in_img_array[27][14][13] <= img[12829];\
        in_img_array[27][14][14] <= img[12830];\
        in_img_array[27][14][15] <= img[12831];\
        in_img_array[27][14][16] <= img[12832];\
        in_img_array[27][14][17] <= img[12833];\
        in_img_array[27][15][0] <= img[12834];\
        in_img_array[27][15][1] <= img[12835];\
        in_img_array[27][15][2] <= img[12836];\
        in_img_array[27][15][3] <= img[12837];\
        in_img_array[27][15][4] <= img[12838];\
        in_img_array[27][15][5] <= img[12839];\
        in_img_array[27][15][6] <= img[12840];\
        in_img_array[27][15][7] <= img[12841];\
        in_img_array[27][15][8] <= img[12842];\
        in_img_array[27][15][9] <= img[12843];\
        in_img_array[27][15][10] <= img[12844];\
        in_img_array[27][15][11] <= img[12845];\
        in_img_array[27][15][12] <= img[12846];\
        in_img_array[27][15][13] <= img[12847];\
        in_img_array[27][15][14] <= img[12848];\
        in_img_array[27][15][15] <= img[12849];\
        in_img_array[27][15][16] <= img[12850];\
        in_img_array[27][15][17] <= img[12851];\
        in_img_array[27][16][0] <= img[12852];\
        in_img_array[27][16][1] <= img[12853];\
        in_img_array[27][16][2] <= img[12854];\
        in_img_array[27][16][3] <= img[12855];\
        in_img_array[27][16][4] <= img[12856];\
        in_img_array[27][16][5] <= img[12857];\
        in_img_array[27][16][6] <= img[12858];\
        in_img_array[27][16][7] <= img[12859];\
        in_img_array[27][16][8] <= img[12860];\
        in_img_array[27][16][9] <= img[12861];\
        in_img_array[27][16][10] <= img[12862];\
        in_img_array[27][16][11] <= img[12863];\
        in_img_array[27][16][12] <= img[12864];\
        in_img_array[27][16][13] <= img[12865];\
        in_img_array[27][16][14] <= img[12866];\
        in_img_array[27][16][15] <= img[12867];\
        in_img_array[27][16][16] <= img[12868];\
        in_img_array[27][16][17] <= img[12869];\
        in_img_array[27][17][0] <= img[12870];\
        in_img_array[27][17][1] <= img[12871];\
        in_img_array[27][17][2] <= img[12872];\
        in_img_array[27][17][3] <= img[12873];\
        in_img_array[27][17][4] <= img[12874];\
        in_img_array[27][17][5] <= img[12875];\
        in_img_array[27][17][6] <= img[12876];\
        in_img_array[27][17][7] <= img[12877];\
        in_img_array[27][17][8] <= img[12878];\
        in_img_array[27][17][9] <= img[12879];\
        in_img_array[27][17][10] <= img[12880];\
        in_img_array[27][17][11] <= img[12881];\
        in_img_array[27][17][12] <= img[12882];\
        in_img_array[27][17][13] <= img[12883];\
        in_img_array[27][17][14] <= img[12884];\
        in_img_array[27][17][15] <= img[12885];\
        in_img_array[27][17][16] <= img[12886];\
        in_img_array[27][17][17] <= img[12887];\
        in_img_array[27][18][0] <= img[12888];\
        in_img_array[27][18][1] <= img[12889];\
        in_img_array[27][18][2] <= img[12890];\
        in_img_array[27][18][3] <= img[12891];\
        in_img_array[27][18][4] <= img[12892];\
        in_img_array[27][18][5] <= img[12893];\
        in_img_array[27][18][6] <= img[12894];\
        in_img_array[27][18][7] <= img[12895];\
        in_img_array[27][18][8] <= img[12896];\
        in_img_array[27][18][9] <= img[12897];\
        in_img_array[27][18][10] <= img[12898];\
        in_img_array[27][18][11] <= img[12899];\
        in_img_array[27][18][12] <= img[12900];\
        in_img_array[27][18][13] <= img[12901];\
        in_img_array[27][18][14] <= img[12902];\
        in_img_array[27][18][15] <= img[12903];\
        in_img_array[27][18][16] <= img[12904];\
        in_img_array[27][18][17] <= img[12905];\
        in_img_array[27][19][0] <= img[12906];\
        in_img_array[27][19][1] <= img[12907];\
        in_img_array[27][19][2] <= img[12908];\
        in_img_array[27][19][3] <= img[12909];\
        in_img_array[27][19][4] <= img[12910];\
        in_img_array[27][19][5] <= img[12911];\
        in_img_array[27][19][6] <= img[12912];\
        in_img_array[27][19][7] <= img[12913];\
        in_img_array[27][19][8] <= img[12914];\
        in_img_array[27][19][9] <= img[12915];\
        in_img_array[27][19][10] <= img[12916];\
        in_img_array[27][19][11] <= img[12917];\
        in_img_array[27][19][12] <= img[12918];\
        in_img_array[27][19][13] <= img[12919];\
        in_img_array[27][19][14] <= img[12920];\
        in_img_array[27][19][15] <= img[12921];\
        in_img_array[27][19][16] <= img[12922];\
        in_img_array[27][19][17] <= img[12923];\
        in_img_array[27][20][0] <= img[12924];\
        in_img_array[27][20][1] <= img[12925];\
        in_img_array[27][20][2] <= img[12926];\
        in_img_array[27][20][3] <= img[12927];\
        in_img_array[27][20][4] <= img[12928];\
        in_img_array[27][20][5] <= img[12929];\
        in_img_array[27][20][6] <= img[12930];\
        in_img_array[27][20][7] <= img[12931];\
        in_img_array[27][20][8] <= img[12932];\
        in_img_array[27][20][9] <= img[12933];\
        in_img_array[27][20][10] <= img[12934];\
        in_img_array[27][20][11] <= img[12935];\
        in_img_array[27][20][12] <= img[12936];\
        in_img_array[27][20][13] <= img[12937];\
        in_img_array[27][20][14] <= img[12938];\
        in_img_array[27][20][15] <= img[12939];\
        in_img_array[27][20][16] <= img[12940];\
        in_img_array[27][20][17] <= img[12941];\
        in_img_array[27][21][0] <= img[12942];\
        in_img_array[27][21][1] <= img[12943];\
        in_img_array[27][21][2] <= img[12944];\
        in_img_array[27][21][3] <= img[12945];\
        in_img_array[27][21][4] <= img[12946];\
        in_img_array[27][21][5] <= img[12947];\
        in_img_array[27][21][6] <= img[12948];\
        in_img_array[27][21][7] <= img[12949];\
        in_img_array[27][21][8] <= img[12950];\
        in_img_array[27][21][9] <= img[12951];\
        in_img_array[27][21][10] <= img[12952];\
        in_img_array[27][21][11] <= img[12953];\
        in_img_array[27][21][12] <= img[12954];\
        in_img_array[27][21][13] <= img[12955];\
        in_img_array[27][21][14] <= img[12956];\
        in_img_array[27][21][15] <= img[12957];\
        in_img_array[27][21][16] <= img[12958];\
        in_img_array[27][21][17] <= img[12959];\
        in_img_array[27][22][0] <= img[12960];\
        in_img_array[27][22][1] <= img[12961];\
        in_img_array[27][22][2] <= img[12962];\
        in_img_array[27][22][3] <= img[12963];\
        in_img_array[27][22][4] <= img[12964];\
        in_img_array[27][22][5] <= img[12965];\
        in_img_array[27][22][6] <= img[12966];\
        in_img_array[27][22][7] <= img[12967];\
        in_img_array[27][22][8] <= img[12968];\
        in_img_array[27][22][9] <= img[12969];\
        in_img_array[27][22][10] <= img[12970];\
        in_img_array[27][22][11] <= img[12971];\
        in_img_array[27][22][12] <= img[12972];\
        in_img_array[27][22][13] <= img[12973];\
        in_img_array[27][22][14] <= img[12974];\
        in_img_array[27][22][15] <= img[12975];\
        in_img_array[27][22][16] <= img[12976];\
        in_img_array[27][22][17] <= img[12977];\
        in_img_array[27][23][0] <= img[12978];\
        in_img_array[27][23][1] <= img[12979];\
        in_img_array[27][23][2] <= img[12980];\
        in_img_array[27][23][3] <= img[12981];\
        in_img_array[27][23][4] <= img[12982];\
        in_img_array[27][23][5] <= img[12983];\
        in_img_array[27][23][6] <= img[12984];\
        in_img_array[27][23][7] <= img[12985];\
        in_img_array[27][23][8] <= img[12986];\
        in_img_array[27][23][9] <= img[12987];\
        in_img_array[27][23][10] <= img[12988];\
        in_img_array[27][23][11] <= img[12989];\
        in_img_array[27][23][12] <= img[12990];\
        in_img_array[27][23][13] <= img[12991];\
        in_img_array[27][23][14] <= img[12992];\
        in_img_array[27][23][15] <= img[12993];\
        in_img_array[27][23][16] <= img[12994];\
        in_img_array[27][23][17] <= img[12995];\
        in_img_array[27][24][0] <= img[12996];\
        in_img_array[27][24][1] <= img[12997];\
        in_img_array[27][24][2] <= img[12998];\
        in_img_array[27][24][3] <= img[12999];\
        in_img_array[27][24][4] <= img[13000];\
        in_img_array[27][24][5] <= img[13001];\
        in_img_array[27][24][6] <= img[13002];\
        in_img_array[27][24][7] <= img[13003];\
        in_img_array[27][24][8] <= img[13004];\
        in_img_array[27][24][9] <= img[13005];\
        in_img_array[27][24][10] <= img[13006];\
        in_img_array[27][24][11] <= img[13007];\
        in_img_array[27][24][12] <= img[13008];\
        in_img_array[27][24][13] <= img[13009];\
        in_img_array[27][24][14] <= img[13010];\
        in_img_array[27][24][15] <= img[13011];\
        in_img_array[27][24][16] <= img[13012];\
        in_img_array[27][24][17] <= img[13013];\
        in_img_array[27][25][0] <= img[13014];\
        in_img_array[27][25][1] <= img[13015];\
        in_img_array[27][25][2] <= img[13016];\
        in_img_array[27][25][3] <= img[13017];\
        in_img_array[27][25][4] <= img[13018];\
        in_img_array[27][25][5] <= img[13019];\
        in_img_array[27][25][6] <= img[13020];\
        in_img_array[27][25][7] <= img[13021];\
        in_img_array[27][25][8] <= img[13022];\
        in_img_array[27][25][9] <= img[13023];\
        in_img_array[27][25][10] <= img[13024];\
        in_img_array[27][25][11] <= img[13025];\
        in_img_array[27][25][12] <= img[13026];\
        in_img_array[27][25][13] <= img[13027];\
        in_img_array[27][25][14] <= img[13028];\
        in_img_array[27][25][15] <= img[13029];\
        in_img_array[27][25][16] <= img[13030];\
        in_img_array[27][25][17] <= img[13031];\
        in_img_array[27][26][0] <= img[13032];\
        in_img_array[27][26][1] <= img[13033];\
        in_img_array[27][26][2] <= img[13034];\
        in_img_array[27][26][3] <= img[13035];\
        in_img_array[27][26][4] <= img[13036];\
        in_img_array[27][26][5] <= img[13037];\
        in_img_array[27][26][6] <= img[13038];\
        in_img_array[27][26][7] <= img[13039];\
        in_img_array[27][26][8] <= img[13040];\
        in_img_array[27][26][9] <= img[13041];\
        in_img_array[27][26][10] <= img[13042];\
        in_img_array[27][26][11] <= img[13043];\
        in_img_array[27][26][12] <= img[13044];\
        in_img_array[27][26][13] <= img[13045];\
        in_img_array[27][26][14] <= img[13046];\
        in_img_array[27][26][15] <= img[13047];\
        in_img_array[27][26][16] <= img[13048];\
        in_img_array[27][26][17] <= img[13049];\
        in_img_array[27][27][0] <= img[13050];\
        in_img_array[27][27][1] <= img[13051];\
        in_img_array[27][27][2] <= img[13052];\
        in_img_array[27][27][3] <= img[13053];\
        in_img_array[27][27][4] <= img[13054];\
        in_img_array[27][27][5] <= img[13055];\
        in_img_array[27][27][6] <= img[13056];\
        in_img_array[27][27][7] <= img[13057];\
        in_img_array[27][27][8] <= img[13058];\
        in_img_array[27][27][9] <= img[13059];\
        in_img_array[27][27][10] <= img[13060];\
        in_img_array[27][27][11] <= img[13061];\
        in_img_array[27][27][12] <= img[13062];\
        in_img_array[27][27][13] <= img[13063];\
        in_img_array[27][27][14] <= img[13064];\
        in_img_array[27][27][15] <= img[13065];\
        in_img_array[27][27][16] <= img[13066];\
        in_img_array[27][27][17] <= img[13067];\
        in_img_array[27][28][0] <= img[13068];\
        in_img_array[27][28][1] <= img[13069];\
        in_img_array[27][28][2] <= img[13070];\
        in_img_array[27][28][3] <= img[13071];\
        in_img_array[27][28][4] <= img[13072];\
        in_img_array[27][28][5] <= img[13073];\
        in_img_array[27][28][6] <= img[13074];\
        in_img_array[27][28][7] <= img[13075];\
        in_img_array[27][28][8] <= img[13076];\
        in_img_array[27][28][9] <= img[13077];\
        in_img_array[27][28][10] <= img[13078];\
        in_img_array[27][28][11] <= img[13079];\
        in_img_array[27][28][12] <= img[13080];\
        in_img_array[27][28][13] <= img[13081];\
        in_img_array[27][28][14] <= img[13082];\
        in_img_array[27][28][15] <= img[13083];\
        in_img_array[27][28][16] <= img[13084];\
        in_img_array[27][28][17] <= img[13085];\
        in_img_array[27][29][0] <= img[13086];\
        in_img_array[27][29][1] <= img[13087];\
        in_img_array[27][29][2] <= img[13088];\
        in_img_array[27][29][3] <= img[13089];\
        in_img_array[27][29][4] <= img[13090];\
        in_img_array[27][29][5] <= img[13091];\
        in_img_array[27][29][6] <= img[13092];\
        in_img_array[27][29][7] <= img[13093];\
        in_img_array[27][29][8] <= img[13094];\
        in_img_array[27][29][9] <= img[13095];\
        in_img_array[27][29][10] <= img[13096];\
        in_img_array[27][29][11] <= img[13097];\
        in_img_array[27][29][12] <= img[13098];\
        in_img_array[27][29][13] <= img[13099];\
        in_img_array[27][29][14] <= img[13100];\
        in_img_array[27][29][15] <= img[13101];\
        in_img_array[27][29][16] <= img[13102];\
        in_img_array[27][29][17] <= img[13103];\
        in_img_array[28][2][0] <= img[13104];\
        in_img_array[28][2][1] <= img[13105];\
        in_img_array[28][2][2] <= img[13106];\
        in_img_array[28][2][3] <= img[13107];\
        in_img_array[28][2][4] <= img[13108];\
        in_img_array[28][2][5] <= img[13109];\
        in_img_array[28][2][6] <= img[13110];\
        in_img_array[28][2][7] <= img[13111];\
        in_img_array[28][2][8] <= img[13112];\
        in_img_array[28][2][9] <= img[13113];\
        in_img_array[28][2][10] <= img[13114];\
        in_img_array[28][2][11] <= img[13115];\
        in_img_array[28][2][12] <= img[13116];\
        in_img_array[28][2][13] <= img[13117];\
        in_img_array[28][2][14] <= img[13118];\
        in_img_array[28][2][15] <= img[13119];\
        in_img_array[28][2][16] <= img[13120];\
        in_img_array[28][2][17] <= img[13121];\
        in_img_array[28][3][0] <= img[13122];\
        in_img_array[28][3][1] <= img[13123];\
        in_img_array[28][3][2] <= img[13124];\
        in_img_array[28][3][3] <= img[13125];\
        in_img_array[28][3][4] <= img[13126];\
        in_img_array[28][3][5] <= img[13127];\
        in_img_array[28][3][6] <= img[13128];\
        in_img_array[28][3][7] <= img[13129];\
        in_img_array[28][3][8] <= img[13130];\
        in_img_array[28][3][9] <= img[13131];\
        in_img_array[28][3][10] <= img[13132];\
        in_img_array[28][3][11] <= img[13133];\
        in_img_array[28][3][12] <= img[13134];\
        in_img_array[28][3][13] <= img[13135];\
        in_img_array[28][3][14] <= img[13136];\
        in_img_array[28][3][15] <= img[13137];\
        in_img_array[28][3][16] <= img[13138];\
        in_img_array[28][3][17] <= img[13139];\
        in_img_array[28][4][0] <= img[13140];\
        in_img_array[28][4][1] <= img[13141];\
        in_img_array[28][4][2] <= img[13142];\
        in_img_array[28][4][3] <= img[13143];\
        in_img_array[28][4][4] <= img[13144];\
        in_img_array[28][4][5] <= img[13145];\
        in_img_array[28][4][6] <= img[13146];\
        in_img_array[28][4][7] <= img[13147];\
        in_img_array[28][4][8] <= img[13148];\
        in_img_array[28][4][9] <= img[13149];\
        in_img_array[28][4][10] <= img[13150];\
        in_img_array[28][4][11] <= img[13151];\
        in_img_array[28][4][12] <= img[13152];\
        in_img_array[28][4][13] <= img[13153];\
        in_img_array[28][4][14] <= img[13154];\
        in_img_array[28][4][15] <= img[13155];\
        in_img_array[28][4][16] <= img[13156];\
        in_img_array[28][4][17] <= img[13157];\
        in_img_array[28][5][0] <= img[13158];\
        in_img_array[28][5][1] <= img[13159];\
        in_img_array[28][5][2] <= img[13160];\
        in_img_array[28][5][3] <= img[13161];\
        in_img_array[28][5][4] <= img[13162];\
        in_img_array[28][5][5] <= img[13163];\
        in_img_array[28][5][6] <= img[13164];\
        in_img_array[28][5][7] <= img[13165];\
        in_img_array[28][5][8] <= img[13166];\
        in_img_array[28][5][9] <= img[13167];\
        in_img_array[28][5][10] <= img[13168];\
        in_img_array[28][5][11] <= img[13169];\
        in_img_array[28][5][12] <= img[13170];\
        in_img_array[28][5][13] <= img[13171];\
        in_img_array[28][5][14] <= img[13172];\
        in_img_array[28][5][15] <= img[13173];\
        in_img_array[28][5][16] <= img[13174];\
        in_img_array[28][5][17] <= img[13175];\
        in_img_array[28][6][0] <= img[13176];\
        in_img_array[28][6][1] <= img[13177];\
        in_img_array[28][6][2] <= img[13178];\
        in_img_array[28][6][3] <= img[13179];\
        in_img_array[28][6][4] <= img[13180];\
        in_img_array[28][6][5] <= img[13181];\
        in_img_array[28][6][6] <= img[13182];\
        in_img_array[28][6][7] <= img[13183];\
        in_img_array[28][6][8] <= img[13184];\
        in_img_array[28][6][9] <= img[13185];\
        in_img_array[28][6][10] <= img[13186];\
        in_img_array[28][6][11] <= img[13187];\
        in_img_array[28][6][12] <= img[13188];\
        in_img_array[28][6][13] <= img[13189];\
        in_img_array[28][6][14] <= img[13190];\
        in_img_array[28][6][15] <= img[13191];\
        in_img_array[28][6][16] <= img[13192];\
        in_img_array[28][6][17] <= img[13193];\
        in_img_array[28][7][0] <= img[13194];\
        in_img_array[28][7][1] <= img[13195];\
        in_img_array[28][7][2] <= img[13196];\
        in_img_array[28][7][3] <= img[13197];\
        in_img_array[28][7][4] <= img[13198];\
        in_img_array[28][7][5] <= img[13199];\
        in_img_array[28][7][6] <= img[13200];\
        in_img_array[28][7][7] <= img[13201];\
        in_img_array[28][7][8] <= img[13202];\
        in_img_array[28][7][9] <= img[13203];\
        in_img_array[28][7][10] <= img[13204];\
        in_img_array[28][7][11] <= img[13205];\
        in_img_array[28][7][12] <= img[13206];\
        in_img_array[28][7][13] <= img[13207];\
        in_img_array[28][7][14] <= img[13208];\
        in_img_array[28][7][15] <= img[13209];\
        in_img_array[28][7][16] <= img[13210];\
        in_img_array[28][7][17] <= img[13211];\
        in_img_array[28][8][0] <= img[13212];\
        in_img_array[28][8][1] <= img[13213];\
        in_img_array[28][8][2] <= img[13214];\
        in_img_array[28][8][3] <= img[13215];\
        in_img_array[28][8][4] <= img[13216];\
        in_img_array[28][8][5] <= img[13217];\
        in_img_array[28][8][6] <= img[13218];\
        in_img_array[28][8][7] <= img[13219];\
        in_img_array[28][8][8] <= img[13220];\
        in_img_array[28][8][9] <= img[13221];\
        in_img_array[28][8][10] <= img[13222];\
        in_img_array[28][8][11] <= img[13223];\
        in_img_array[28][8][12] <= img[13224];\
        in_img_array[28][8][13] <= img[13225];\
        in_img_array[28][8][14] <= img[13226];\
        in_img_array[28][8][15] <= img[13227];\
        in_img_array[28][8][16] <= img[13228];\
        in_img_array[28][8][17] <= img[13229];\
        in_img_array[28][9][0] <= img[13230];\
        in_img_array[28][9][1] <= img[13231];\
        in_img_array[28][9][2] <= img[13232];\
        in_img_array[28][9][3] <= img[13233];\
        in_img_array[28][9][4] <= img[13234];\
        in_img_array[28][9][5] <= img[13235];\
        in_img_array[28][9][6] <= img[13236];\
        in_img_array[28][9][7] <= img[13237];\
        in_img_array[28][9][8] <= img[13238];\
        in_img_array[28][9][9] <= img[13239];\
        in_img_array[28][9][10] <= img[13240];\
        in_img_array[28][9][11] <= img[13241];\
        in_img_array[28][9][12] <= img[13242];\
        in_img_array[28][9][13] <= img[13243];\
        in_img_array[28][9][14] <= img[13244];\
        in_img_array[28][9][15] <= img[13245];\
        in_img_array[28][9][16] <= img[13246];\
        in_img_array[28][9][17] <= img[13247];\
        in_img_array[28][10][0] <= img[13248];\
        in_img_array[28][10][1] <= img[13249];\
        in_img_array[28][10][2] <= img[13250];\
        in_img_array[28][10][3] <= img[13251];\
        in_img_array[28][10][4] <= img[13252];\
        in_img_array[28][10][5] <= img[13253];\
        in_img_array[28][10][6] <= img[13254];\
        in_img_array[28][10][7] <= img[13255];\
        in_img_array[28][10][8] <= img[13256];\
        in_img_array[28][10][9] <= img[13257];\
        in_img_array[28][10][10] <= img[13258];\
        in_img_array[28][10][11] <= img[13259];\
        in_img_array[28][10][12] <= img[13260];\
        in_img_array[28][10][13] <= img[13261];\
        in_img_array[28][10][14] <= img[13262];\
        in_img_array[28][10][15] <= img[13263];\
        in_img_array[28][10][16] <= img[13264];\
        in_img_array[28][10][17] <= img[13265];\
        in_img_array[28][11][0] <= img[13266];\
        in_img_array[28][11][1] <= img[13267];\
        in_img_array[28][11][2] <= img[13268];\
        in_img_array[28][11][3] <= img[13269];\
        in_img_array[28][11][4] <= img[13270];\
        in_img_array[28][11][5] <= img[13271];\
        in_img_array[28][11][6] <= img[13272];\
        in_img_array[28][11][7] <= img[13273];\
        in_img_array[28][11][8] <= img[13274];\
        in_img_array[28][11][9] <= img[13275];\
        in_img_array[28][11][10] <= img[13276];\
        in_img_array[28][11][11] <= img[13277];\
        in_img_array[28][11][12] <= img[13278];\
        in_img_array[28][11][13] <= img[13279];\
        in_img_array[28][11][14] <= img[13280];\
        in_img_array[28][11][15] <= img[13281];\
        in_img_array[28][11][16] <= img[13282];\
        in_img_array[28][11][17] <= img[13283];\
        in_img_array[28][12][0] <= img[13284];\
        in_img_array[28][12][1] <= img[13285];\
        in_img_array[28][12][2] <= img[13286];\
        in_img_array[28][12][3] <= img[13287];\
        in_img_array[28][12][4] <= img[13288];\
        in_img_array[28][12][5] <= img[13289];\
        in_img_array[28][12][6] <= img[13290];\
        in_img_array[28][12][7] <= img[13291];\
        in_img_array[28][12][8] <= img[13292];\
        in_img_array[28][12][9] <= img[13293];\
        in_img_array[28][12][10] <= img[13294];\
        in_img_array[28][12][11] <= img[13295];\
        in_img_array[28][12][12] <= img[13296];\
        in_img_array[28][12][13] <= img[13297];\
        in_img_array[28][12][14] <= img[13298];\
        in_img_array[28][12][15] <= img[13299];\
        in_img_array[28][12][16] <= img[13300];\
        in_img_array[28][12][17] <= img[13301];\
        in_img_array[28][13][0] <= img[13302];\
        in_img_array[28][13][1] <= img[13303];\
        in_img_array[28][13][2] <= img[13304];\
        in_img_array[28][13][3] <= img[13305];\
        in_img_array[28][13][4] <= img[13306];\
        in_img_array[28][13][5] <= img[13307];\
        in_img_array[28][13][6] <= img[13308];\
        in_img_array[28][13][7] <= img[13309];\
        in_img_array[28][13][8] <= img[13310];\
        in_img_array[28][13][9] <= img[13311];\
        in_img_array[28][13][10] <= img[13312];\
        in_img_array[28][13][11] <= img[13313];\
        in_img_array[28][13][12] <= img[13314];\
        in_img_array[28][13][13] <= img[13315];\
        in_img_array[28][13][14] <= img[13316];\
        in_img_array[28][13][15] <= img[13317];\
        in_img_array[28][13][16] <= img[13318];\
        in_img_array[28][13][17] <= img[13319];\
        in_img_array[28][14][0] <= img[13320];\
        in_img_array[28][14][1] <= img[13321];\
        in_img_array[28][14][2] <= img[13322];\
        in_img_array[28][14][3] <= img[13323];\
        in_img_array[28][14][4] <= img[13324];\
        in_img_array[28][14][5] <= img[13325];\
        in_img_array[28][14][6] <= img[13326];\
        in_img_array[28][14][7] <= img[13327];\
        in_img_array[28][14][8] <= img[13328];\
        in_img_array[28][14][9] <= img[13329];\
        in_img_array[28][14][10] <= img[13330];\
        in_img_array[28][14][11] <= img[13331];\
        in_img_array[28][14][12] <= img[13332];\
        in_img_array[28][14][13] <= img[13333];\
        in_img_array[28][14][14] <= img[13334];\
        in_img_array[28][14][15] <= img[13335];\
        in_img_array[28][14][16] <= img[13336];\
        in_img_array[28][14][17] <= img[13337];\
        in_img_array[28][15][0] <= img[13338];\
        in_img_array[28][15][1] <= img[13339];\
        in_img_array[28][15][2] <= img[13340];\
        in_img_array[28][15][3] <= img[13341];\
        in_img_array[28][15][4] <= img[13342];\
        in_img_array[28][15][5] <= img[13343];\
        in_img_array[28][15][6] <= img[13344];\
        in_img_array[28][15][7] <= img[13345];\
        in_img_array[28][15][8] <= img[13346];\
        in_img_array[28][15][9] <= img[13347];\
        in_img_array[28][15][10] <= img[13348];\
        in_img_array[28][15][11] <= img[13349];\
        in_img_array[28][15][12] <= img[13350];\
        in_img_array[28][15][13] <= img[13351];\
        in_img_array[28][15][14] <= img[13352];\
        in_img_array[28][15][15] <= img[13353];\
        in_img_array[28][15][16] <= img[13354];\
        in_img_array[28][15][17] <= img[13355];\
        in_img_array[28][16][0] <= img[13356];\
        in_img_array[28][16][1] <= img[13357];\
        in_img_array[28][16][2] <= img[13358];\
        in_img_array[28][16][3] <= img[13359];\
        in_img_array[28][16][4] <= img[13360];\
        in_img_array[28][16][5] <= img[13361];\
        in_img_array[28][16][6] <= img[13362];\
        in_img_array[28][16][7] <= img[13363];\
        in_img_array[28][16][8] <= img[13364];\
        in_img_array[28][16][9] <= img[13365];\
        in_img_array[28][16][10] <= img[13366];\
        in_img_array[28][16][11] <= img[13367];\
        in_img_array[28][16][12] <= img[13368];\
        in_img_array[28][16][13] <= img[13369];\
        in_img_array[28][16][14] <= img[13370];\
        in_img_array[28][16][15] <= img[13371];\
        in_img_array[28][16][16] <= img[13372];\
        in_img_array[28][16][17] <= img[13373];\
        in_img_array[28][17][0] <= img[13374];\
        in_img_array[28][17][1] <= img[13375];\
        in_img_array[28][17][2] <= img[13376];\
        in_img_array[28][17][3] <= img[13377];\
        in_img_array[28][17][4] <= img[13378];\
        in_img_array[28][17][5] <= img[13379];\
        in_img_array[28][17][6] <= img[13380];\
        in_img_array[28][17][7] <= img[13381];\
        in_img_array[28][17][8] <= img[13382];\
        in_img_array[28][17][9] <= img[13383];\
        in_img_array[28][17][10] <= img[13384];\
        in_img_array[28][17][11] <= img[13385];\
        in_img_array[28][17][12] <= img[13386];\
        in_img_array[28][17][13] <= img[13387];\
        in_img_array[28][17][14] <= img[13388];\
        in_img_array[28][17][15] <= img[13389];\
        in_img_array[28][17][16] <= img[13390];\
        in_img_array[28][17][17] <= img[13391];\
        in_img_array[28][18][0] <= img[13392];\
        in_img_array[28][18][1] <= img[13393];\
        in_img_array[28][18][2] <= img[13394];\
        in_img_array[28][18][3] <= img[13395];\
        in_img_array[28][18][4] <= img[13396];\
        in_img_array[28][18][5] <= img[13397];\
        in_img_array[28][18][6] <= img[13398];\
        in_img_array[28][18][7] <= img[13399];\
        in_img_array[28][18][8] <= img[13400];\
        in_img_array[28][18][9] <= img[13401];\
        in_img_array[28][18][10] <= img[13402];\
        in_img_array[28][18][11] <= img[13403];\
        in_img_array[28][18][12] <= img[13404];\
        in_img_array[28][18][13] <= img[13405];\
        in_img_array[28][18][14] <= img[13406];\
        in_img_array[28][18][15] <= img[13407];\
        in_img_array[28][18][16] <= img[13408];\
        in_img_array[28][18][17] <= img[13409];\
        in_img_array[28][19][0] <= img[13410];\
        in_img_array[28][19][1] <= img[13411];\
        in_img_array[28][19][2] <= img[13412];\
        in_img_array[28][19][3] <= img[13413];\
        in_img_array[28][19][4] <= img[13414];\
        in_img_array[28][19][5] <= img[13415];\
        in_img_array[28][19][6] <= img[13416];\
        in_img_array[28][19][7] <= img[13417];\
        in_img_array[28][19][8] <= img[13418];\
        in_img_array[28][19][9] <= img[13419];\
        in_img_array[28][19][10] <= img[13420];\
        in_img_array[28][19][11] <= img[13421];\
        in_img_array[28][19][12] <= img[13422];\
        in_img_array[28][19][13] <= img[13423];\
        in_img_array[28][19][14] <= img[13424];\
        in_img_array[28][19][15] <= img[13425];\
        in_img_array[28][19][16] <= img[13426];\
        in_img_array[28][19][17] <= img[13427];\
        in_img_array[28][20][0] <= img[13428];\
        in_img_array[28][20][1] <= img[13429];\
        in_img_array[28][20][2] <= img[13430];\
        in_img_array[28][20][3] <= img[13431];\
        in_img_array[28][20][4] <= img[13432];\
        in_img_array[28][20][5] <= img[13433];\
        in_img_array[28][20][6] <= img[13434];\
        in_img_array[28][20][7] <= img[13435];\
        in_img_array[28][20][8] <= img[13436];\
        in_img_array[28][20][9] <= img[13437];\
        in_img_array[28][20][10] <= img[13438];\
        in_img_array[28][20][11] <= img[13439];\
        in_img_array[28][20][12] <= img[13440];\
        in_img_array[28][20][13] <= img[13441];\
        in_img_array[28][20][14] <= img[13442];\
        in_img_array[28][20][15] <= img[13443];\
        in_img_array[28][20][16] <= img[13444];\
        in_img_array[28][20][17] <= img[13445];\
        in_img_array[28][21][0] <= img[13446];\
        in_img_array[28][21][1] <= img[13447];\
        in_img_array[28][21][2] <= img[13448];\
        in_img_array[28][21][3] <= img[13449];\
        in_img_array[28][21][4] <= img[13450];\
        in_img_array[28][21][5] <= img[13451];\
        in_img_array[28][21][6] <= img[13452];\
        in_img_array[28][21][7] <= img[13453];\
        in_img_array[28][21][8] <= img[13454];\
        in_img_array[28][21][9] <= img[13455];\
        in_img_array[28][21][10] <= img[13456];\
        in_img_array[28][21][11] <= img[13457];\
        in_img_array[28][21][12] <= img[13458];\
        in_img_array[28][21][13] <= img[13459];\
        in_img_array[28][21][14] <= img[13460];\
        in_img_array[28][21][15] <= img[13461];\
        in_img_array[28][21][16] <= img[13462];\
        in_img_array[28][21][17] <= img[13463];\
        in_img_array[28][22][0] <= img[13464];\
        in_img_array[28][22][1] <= img[13465];\
        in_img_array[28][22][2] <= img[13466];\
        in_img_array[28][22][3] <= img[13467];\
        in_img_array[28][22][4] <= img[13468];\
        in_img_array[28][22][5] <= img[13469];\
        in_img_array[28][22][6] <= img[13470];\
        in_img_array[28][22][7] <= img[13471];\
        in_img_array[28][22][8] <= img[13472];\
        in_img_array[28][22][9] <= img[13473];\
        in_img_array[28][22][10] <= img[13474];\
        in_img_array[28][22][11] <= img[13475];\
        in_img_array[28][22][12] <= img[13476];\
        in_img_array[28][22][13] <= img[13477];\
        in_img_array[28][22][14] <= img[13478];\
        in_img_array[28][22][15] <= img[13479];\
        in_img_array[28][22][16] <= img[13480];\
        in_img_array[28][22][17] <= img[13481];\
        in_img_array[28][23][0] <= img[13482];\
        in_img_array[28][23][1] <= img[13483];\
        in_img_array[28][23][2] <= img[13484];\
        in_img_array[28][23][3] <= img[13485];\
        in_img_array[28][23][4] <= img[13486];\
        in_img_array[28][23][5] <= img[13487];\
        in_img_array[28][23][6] <= img[13488];\
        in_img_array[28][23][7] <= img[13489];\
        in_img_array[28][23][8] <= img[13490];\
        in_img_array[28][23][9] <= img[13491];\
        in_img_array[28][23][10] <= img[13492];\
        in_img_array[28][23][11] <= img[13493];\
        in_img_array[28][23][12] <= img[13494];\
        in_img_array[28][23][13] <= img[13495];\
        in_img_array[28][23][14] <= img[13496];\
        in_img_array[28][23][15] <= img[13497];\
        in_img_array[28][23][16] <= img[13498];\
        in_img_array[28][23][17] <= img[13499];\
        in_img_array[28][24][0] <= img[13500];\
        in_img_array[28][24][1] <= img[13501];\
        in_img_array[28][24][2] <= img[13502];\
        in_img_array[28][24][3] <= img[13503];\
        in_img_array[28][24][4] <= img[13504];\
        in_img_array[28][24][5] <= img[13505];\
        in_img_array[28][24][6] <= img[13506];\
        in_img_array[28][24][7] <= img[13507];\
        in_img_array[28][24][8] <= img[13508];\
        in_img_array[28][24][9] <= img[13509];\
        in_img_array[28][24][10] <= img[13510];\
        in_img_array[28][24][11] <= img[13511];\
        in_img_array[28][24][12] <= img[13512];\
        in_img_array[28][24][13] <= img[13513];\
        in_img_array[28][24][14] <= img[13514];\
        in_img_array[28][24][15] <= img[13515];\
        in_img_array[28][24][16] <= img[13516];\
        in_img_array[28][24][17] <= img[13517];\
        in_img_array[28][25][0] <= img[13518];\
        in_img_array[28][25][1] <= img[13519];\
        in_img_array[28][25][2] <= img[13520];\
        in_img_array[28][25][3] <= img[13521];\
        in_img_array[28][25][4] <= img[13522];\
        in_img_array[28][25][5] <= img[13523];\
        in_img_array[28][25][6] <= img[13524];\
        in_img_array[28][25][7] <= img[13525];\
        in_img_array[28][25][8] <= img[13526];\
        in_img_array[28][25][9] <= img[13527];\
        in_img_array[28][25][10] <= img[13528];\
        in_img_array[28][25][11] <= img[13529];\
        in_img_array[28][25][12] <= img[13530];\
        in_img_array[28][25][13] <= img[13531];\
        in_img_array[28][25][14] <= img[13532];\
        in_img_array[28][25][15] <= img[13533];\
        in_img_array[28][25][16] <= img[13534];\
        in_img_array[28][25][17] <= img[13535];\
        in_img_array[28][26][0] <= img[13536];\
        in_img_array[28][26][1] <= img[13537];\
        in_img_array[28][26][2] <= img[13538];\
        in_img_array[28][26][3] <= img[13539];\
        in_img_array[28][26][4] <= img[13540];\
        in_img_array[28][26][5] <= img[13541];\
        in_img_array[28][26][6] <= img[13542];\
        in_img_array[28][26][7] <= img[13543];\
        in_img_array[28][26][8] <= img[13544];\
        in_img_array[28][26][9] <= img[13545];\
        in_img_array[28][26][10] <= img[13546];\
        in_img_array[28][26][11] <= img[13547];\
        in_img_array[28][26][12] <= img[13548];\
        in_img_array[28][26][13] <= img[13549];\
        in_img_array[28][26][14] <= img[13550];\
        in_img_array[28][26][15] <= img[13551];\
        in_img_array[28][26][16] <= img[13552];\
        in_img_array[28][26][17] <= img[13553];\
        in_img_array[28][27][0] <= img[13554];\
        in_img_array[28][27][1] <= img[13555];\
        in_img_array[28][27][2] <= img[13556];\
        in_img_array[28][27][3] <= img[13557];\
        in_img_array[28][27][4] <= img[13558];\
        in_img_array[28][27][5] <= img[13559];\
        in_img_array[28][27][6] <= img[13560];\
        in_img_array[28][27][7] <= img[13561];\
        in_img_array[28][27][8] <= img[13562];\
        in_img_array[28][27][9] <= img[13563];\
        in_img_array[28][27][10] <= img[13564];\
        in_img_array[28][27][11] <= img[13565];\
        in_img_array[28][27][12] <= img[13566];\
        in_img_array[28][27][13] <= img[13567];\
        in_img_array[28][27][14] <= img[13568];\
        in_img_array[28][27][15] <= img[13569];\
        in_img_array[28][27][16] <= img[13570];\
        in_img_array[28][27][17] <= img[13571];\
        in_img_array[28][28][0] <= img[13572];\
        in_img_array[28][28][1] <= img[13573];\
        in_img_array[28][28][2] <= img[13574];\
        in_img_array[28][28][3] <= img[13575];\
        in_img_array[28][28][4] <= img[13576];\
        in_img_array[28][28][5] <= img[13577];\
        in_img_array[28][28][6] <= img[13578];\
        in_img_array[28][28][7] <= img[13579];\
        in_img_array[28][28][8] <= img[13580];\
        in_img_array[28][28][9] <= img[13581];\
        in_img_array[28][28][10] <= img[13582];\
        in_img_array[28][28][11] <= img[13583];\
        in_img_array[28][28][12] <= img[13584];\
        in_img_array[28][28][13] <= img[13585];\
        in_img_array[28][28][14] <= img[13586];\
        in_img_array[28][28][15] <= img[13587];\
        in_img_array[28][28][16] <= img[13588];\
        in_img_array[28][28][17] <= img[13589];\
        in_img_array[28][29][0] <= img[13590];\
        in_img_array[28][29][1] <= img[13591];\
        in_img_array[28][29][2] <= img[13592];\
        in_img_array[28][29][3] <= img[13593];\
        in_img_array[28][29][4] <= img[13594];\
        in_img_array[28][29][5] <= img[13595];\
        in_img_array[28][29][6] <= img[13596];\
        in_img_array[28][29][7] <= img[13597];\
        in_img_array[28][29][8] <= img[13598];\
        in_img_array[28][29][9] <= img[13599];\
        in_img_array[28][29][10] <= img[13600];\
        in_img_array[28][29][11] <= img[13601];\
        in_img_array[28][29][12] <= img[13602];\
        in_img_array[28][29][13] <= img[13603];\
        in_img_array[28][29][14] <= img[13604];\
        in_img_array[28][29][15] <= img[13605];\
        in_img_array[28][29][16] <= img[13606];\
        in_img_array[28][29][17] <= img[13607];\
        in_img_array[29][2][0] <= img[13608];\
        in_img_array[29][2][1] <= img[13609];\
        in_img_array[29][2][2] <= img[13610];\
        in_img_array[29][2][3] <= img[13611];\
        in_img_array[29][2][4] <= img[13612];\
        in_img_array[29][2][5] <= img[13613];\
        in_img_array[29][2][6] <= img[13614];\
        in_img_array[29][2][7] <= img[13615];\
        in_img_array[29][2][8] <= img[13616];\
        in_img_array[29][2][9] <= img[13617];\
        in_img_array[29][2][10] <= img[13618];\
        in_img_array[29][2][11] <= img[13619];\
        in_img_array[29][2][12] <= img[13620];\
        in_img_array[29][2][13] <= img[13621];\
        in_img_array[29][2][14] <= img[13622];\
        in_img_array[29][2][15] <= img[13623];\
        in_img_array[29][2][16] <= img[13624];\
        in_img_array[29][2][17] <= img[13625];\
        in_img_array[29][3][0] <= img[13626];\
        in_img_array[29][3][1] <= img[13627];\
        in_img_array[29][3][2] <= img[13628];\
        in_img_array[29][3][3] <= img[13629];\
        in_img_array[29][3][4] <= img[13630];\
        in_img_array[29][3][5] <= img[13631];\
        in_img_array[29][3][6] <= img[13632];\
        in_img_array[29][3][7] <= img[13633];\
        in_img_array[29][3][8] <= img[13634];\
        in_img_array[29][3][9] <= img[13635];\
        in_img_array[29][3][10] <= img[13636];\
        in_img_array[29][3][11] <= img[13637];\
        in_img_array[29][3][12] <= img[13638];\
        in_img_array[29][3][13] <= img[13639];\
        in_img_array[29][3][14] <= img[13640];\
        in_img_array[29][3][15] <= img[13641];\
        in_img_array[29][3][16] <= img[13642];\
        in_img_array[29][3][17] <= img[13643];\
        in_img_array[29][4][0] <= img[13644];\
        in_img_array[29][4][1] <= img[13645];\
        in_img_array[29][4][2] <= img[13646];\
        in_img_array[29][4][3] <= img[13647];\
        in_img_array[29][4][4] <= img[13648];\
        in_img_array[29][4][5] <= img[13649];\
        in_img_array[29][4][6] <= img[13650];\
        in_img_array[29][4][7] <= img[13651];\
        in_img_array[29][4][8] <= img[13652];\
        in_img_array[29][4][9] <= img[13653];\
        in_img_array[29][4][10] <= img[13654];\
        in_img_array[29][4][11] <= img[13655];\
        in_img_array[29][4][12] <= img[13656];\
        in_img_array[29][4][13] <= img[13657];\
        in_img_array[29][4][14] <= img[13658];\
        in_img_array[29][4][15] <= img[13659];\
        in_img_array[29][4][16] <= img[13660];\
        in_img_array[29][4][17] <= img[13661];\
        in_img_array[29][5][0] <= img[13662];\
        in_img_array[29][5][1] <= img[13663];\
        in_img_array[29][5][2] <= img[13664];\
        in_img_array[29][5][3] <= img[13665];\
        in_img_array[29][5][4] <= img[13666];\
        in_img_array[29][5][5] <= img[13667];\
        in_img_array[29][5][6] <= img[13668];\
        in_img_array[29][5][7] <= img[13669];\
        in_img_array[29][5][8] <= img[13670];\
        in_img_array[29][5][9] <= img[13671];\
        in_img_array[29][5][10] <= img[13672];\
        in_img_array[29][5][11] <= img[13673];\
        in_img_array[29][5][12] <= img[13674];\
        in_img_array[29][5][13] <= img[13675];\
        in_img_array[29][5][14] <= img[13676];\
        in_img_array[29][5][15] <= img[13677];\
        in_img_array[29][5][16] <= img[13678];\
        in_img_array[29][5][17] <= img[13679];\
        in_img_array[29][6][0] <= img[13680];\
        in_img_array[29][6][1] <= img[13681];\
        in_img_array[29][6][2] <= img[13682];\
        in_img_array[29][6][3] <= img[13683];\
        in_img_array[29][6][4] <= img[13684];\
        in_img_array[29][6][5] <= img[13685];\
        in_img_array[29][6][6] <= img[13686];\
        in_img_array[29][6][7] <= img[13687];\
        in_img_array[29][6][8] <= img[13688];\
        in_img_array[29][6][9] <= img[13689];\
        in_img_array[29][6][10] <= img[13690];\
        in_img_array[29][6][11] <= img[13691];\
        in_img_array[29][6][12] <= img[13692];\
        in_img_array[29][6][13] <= img[13693];\
        in_img_array[29][6][14] <= img[13694];\
        in_img_array[29][6][15] <= img[13695];\
        in_img_array[29][6][16] <= img[13696];\
        in_img_array[29][6][17] <= img[13697];\
        in_img_array[29][7][0] <= img[13698];\
        in_img_array[29][7][1] <= img[13699];\
        in_img_array[29][7][2] <= img[13700];\
        in_img_array[29][7][3] <= img[13701];\
        in_img_array[29][7][4] <= img[13702];\
        in_img_array[29][7][5] <= img[13703];\
        in_img_array[29][7][6] <= img[13704];\
        in_img_array[29][7][7] <= img[13705];\
        in_img_array[29][7][8] <= img[13706];\
        in_img_array[29][7][9] <= img[13707];\
        in_img_array[29][7][10] <= img[13708];\
        in_img_array[29][7][11] <= img[13709];\
        in_img_array[29][7][12] <= img[13710];\
        in_img_array[29][7][13] <= img[13711];\
        in_img_array[29][7][14] <= img[13712];\
        in_img_array[29][7][15] <= img[13713];\
        in_img_array[29][7][16] <= img[13714];\
        in_img_array[29][7][17] <= img[13715];\
        in_img_array[29][8][0] <= img[13716];\
        in_img_array[29][8][1] <= img[13717];\
        in_img_array[29][8][2] <= img[13718];\
        in_img_array[29][8][3] <= img[13719];\
        in_img_array[29][8][4] <= img[13720];\
        in_img_array[29][8][5] <= img[13721];\
        in_img_array[29][8][6] <= img[13722];\
        in_img_array[29][8][7] <= img[13723];\
        in_img_array[29][8][8] <= img[13724];\
        in_img_array[29][8][9] <= img[13725];\
        in_img_array[29][8][10] <= img[13726];\
        in_img_array[29][8][11] <= img[13727];\
        in_img_array[29][8][12] <= img[13728];\
        in_img_array[29][8][13] <= img[13729];\
        in_img_array[29][8][14] <= img[13730];\
        in_img_array[29][8][15] <= img[13731];\
        in_img_array[29][8][16] <= img[13732];\
        in_img_array[29][8][17] <= img[13733];\
        in_img_array[29][9][0] <= img[13734];\
        in_img_array[29][9][1] <= img[13735];\
        in_img_array[29][9][2] <= img[13736];\
        in_img_array[29][9][3] <= img[13737];\
        in_img_array[29][9][4] <= img[13738];\
        in_img_array[29][9][5] <= img[13739];\
        in_img_array[29][9][6] <= img[13740];\
        in_img_array[29][9][7] <= img[13741];\
        in_img_array[29][9][8] <= img[13742];\
        in_img_array[29][9][9] <= img[13743];\
        in_img_array[29][9][10] <= img[13744];\
        in_img_array[29][9][11] <= img[13745];\
        in_img_array[29][9][12] <= img[13746];\
        in_img_array[29][9][13] <= img[13747];\
        in_img_array[29][9][14] <= img[13748];\
        in_img_array[29][9][15] <= img[13749];\
        in_img_array[29][9][16] <= img[13750];\
        in_img_array[29][9][17] <= img[13751];\
        in_img_array[29][10][0] <= img[13752];\
        in_img_array[29][10][1] <= img[13753];\
        in_img_array[29][10][2] <= img[13754];\
        in_img_array[29][10][3] <= img[13755];\
        in_img_array[29][10][4] <= img[13756];\
        in_img_array[29][10][5] <= img[13757];\
        in_img_array[29][10][6] <= img[13758];\
        in_img_array[29][10][7] <= img[13759];\
        in_img_array[29][10][8] <= img[13760];\
        in_img_array[29][10][9] <= img[13761];\
        in_img_array[29][10][10] <= img[13762];\
        in_img_array[29][10][11] <= img[13763];\
        in_img_array[29][10][12] <= img[13764];\
        in_img_array[29][10][13] <= img[13765];\
        in_img_array[29][10][14] <= img[13766];\
        in_img_array[29][10][15] <= img[13767];\
        in_img_array[29][10][16] <= img[13768];\
        in_img_array[29][10][17] <= img[13769];\
        in_img_array[29][11][0] <= img[13770];\
        in_img_array[29][11][1] <= img[13771];\
        in_img_array[29][11][2] <= img[13772];\
        in_img_array[29][11][3] <= img[13773];\
        in_img_array[29][11][4] <= img[13774];\
        in_img_array[29][11][5] <= img[13775];\
        in_img_array[29][11][6] <= img[13776];\
        in_img_array[29][11][7] <= img[13777];\
        in_img_array[29][11][8] <= img[13778];\
        in_img_array[29][11][9] <= img[13779];\
        in_img_array[29][11][10] <= img[13780];\
        in_img_array[29][11][11] <= img[13781];\
        in_img_array[29][11][12] <= img[13782];\
        in_img_array[29][11][13] <= img[13783];\
        in_img_array[29][11][14] <= img[13784];\
        in_img_array[29][11][15] <= img[13785];\
        in_img_array[29][11][16] <= img[13786];\
        in_img_array[29][11][17] <= img[13787];\
        in_img_array[29][12][0] <= img[13788];\
        in_img_array[29][12][1] <= img[13789];\
        in_img_array[29][12][2] <= img[13790];\
        in_img_array[29][12][3] <= img[13791];\
        in_img_array[29][12][4] <= img[13792];\
        in_img_array[29][12][5] <= img[13793];\
        in_img_array[29][12][6] <= img[13794];\
        in_img_array[29][12][7] <= img[13795];\
        in_img_array[29][12][8] <= img[13796];\
        in_img_array[29][12][9] <= img[13797];\
        in_img_array[29][12][10] <= img[13798];\
        in_img_array[29][12][11] <= img[13799];\
        in_img_array[29][12][12] <= img[13800];\
        in_img_array[29][12][13] <= img[13801];\
        in_img_array[29][12][14] <= img[13802];\
        in_img_array[29][12][15] <= img[13803];\
        in_img_array[29][12][16] <= img[13804];\
        in_img_array[29][12][17] <= img[13805];\
        in_img_array[29][13][0] <= img[13806];\
        in_img_array[29][13][1] <= img[13807];\
        in_img_array[29][13][2] <= img[13808];\
        in_img_array[29][13][3] <= img[13809];\
        in_img_array[29][13][4] <= img[13810];\
        in_img_array[29][13][5] <= img[13811];\
        in_img_array[29][13][6] <= img[13812];\
        in_img_array[29][13][7] <= img[13813];\
        in_img_array[29][13][8] <= img[13814];\
        in_img_array[29][13][9] <= img[13815];\
        in_img_array[29][13][10] <= img[13816];\
        in_img_array[29][13][11] <= img[13817];\
        in_img_array[29][13][12] <= img[13818];\
        in_img_array[29][13][13] <= img[13819];\
        in_img_array[29][13][14] <= img[13820];\
        in_img_array[29][13][15] <= img[13821];\
        in_img_array[29][13][16] <= img[13822];\
        in_img_array[29][13][17] <= img[13823];\
        in_img_array[29][14][0] <= img[13824];\
        in_img_array[29][14][1] <= img[13825];\
        in_img_array[29][14][2] <= img[13826];\
        in_img_array[29][14][3] <= img[13827];\
        in_img_array[29][14][4] <= img[13828];\
        in_img_array[29][14][5] <= img[13829];\
        in_img_array[29][14][6] <= img[13830];\
        in_img_array[29][14][7] <= img[13831];\
        in_img_array[29][14][8] <= img[13832];\
        in_img_array[29][14][9] <= img[13833];\
        in_img_array[29][14][10] <= img[13834];\
        in_img_array[29][14][11] <= img[13835];\
        in_img_array[29][14][12] <= img[13836];\
        in_img_array[29][14][13] <= img[13837];\
        in_img_array[29][14][14] <= img[13838];\
        in_img_array[29][14][15] <= img[13839];\
        in_img_array[29][14][16] <= img[13840];\
        in_img_array[29][14][17] <= img[13841];\
        in_img_array[29][15][0] <= img[13842];\
        in_img_array[29][15][1] <= img[13843];\
        in_img_array[29][15][2] <= img[13844];\
        in_img_array[29][15][3] <= img[13845];\
        in_img_array[29][15][4] <= img[13846];\
        in_img_array[29][15][5] <= img[13847];\
        in_img_array[29][15][6] <= img[13848];\
        in_img_array[29][15][7] <= img[13849];\
        in_img_array[29][15][8] <= img[13850];\
        in_img_array[29][15][9] <= img[13851];\
        in_img_array[29][15][10] <= img[13852];\
        in_img_array[29][15][11] <= img[13853];\
        in_img_array[29][15][12] <= img[13854];\
        in_img_array[29][15][13] <= img[13855];\
        in_img_array[29][15][14] <= img[13856];\
        in_img_array[29][15][15] <= img[13857];\
        in_img_array[29][15][16] <= img[13858];\
        in_img_array[29][15][17] <= img[13859];\
        in_img_array[29][16][0] <= img[13860];\
        in_img_array[29][16][1] <= img[13861];\
        in_img_array[29][16][2] <= img[13862];\
        in_img_array[29][16][3] <= img[13863];\
        in_img_array[29][16][4] <= img[13864];\
        in_img_array[29][16][5] <= img[13865];\
        in_img_array[29][16][6] <= img[13866];\
        in_img_array[29][16][7] <= img[13867];\
        in_img_array[29][16][8] <= img[13868];\
        in_img_array[29][16][9] <= img[13869];\
        in_img_array[29][16][10] <= img[13870];\
        in_img_array[29][16][11] <= img[13871];\
        in_img_array[29][16][12] <= img[13872];\
        in_img_array[29][16][13] <= img[13873];\
        in_img_array[29][16][14] <= img[13874];\
        in_img_array[29][16][15] <= img[13875];\
        in_img_array[29][16][16] <= img[13876];\
        in_img_array[29][16][17] <= img[13877];\
        in_img_array[29][17][0] <= img[13878];\
        in_img_array[29][17][1] <= img[13879];\
        in_img_array[29][17][2] <= img[13880];\
        in_img_array[29][17][3] <= img[13881];\
        in_img_array[29][17][4] <= img[13882];\
        in_img_array[29][17][5] <= img[13883];\
        in_img_array[29][17][6] <= img[13884];\
        in_img_array[29][17][7] <= img[13885];\
        in_img_array[29][17][8] <= img[13886];\
        in_img_array[29][17][9] <= img[13887];\
        in_img_array[29][17][10] <= img[13888];\
        in_img_array[29][17][11] <= img[13889];\
        in_img_array[29][17][12] <= img[13890];\
        in_img_array[29][17][13] <= img[13891];\
        in_img_array[29][17][14] <= img[13892];\
        in_img_array[29][17][15] <= img[13893];\
        in_img_array[29][17][16] <= img[13894];\
        in_img_array[29][17][17] <= img[13895];\
        in_img_array[29][18][0] <= img[13896];\
        in_img_array[29][18][1] <= img[13897];\
        in_img_array[29][18][2] <= img[13898];\
        in_img_array[29][18][3] <= img[13899];\
        in_img_array[29][18][4] <= img[13900];\
        in_img_array[29][18][5] <= img[13901];\
        in_img_array[29][18][6] <= img[13902];\
        in_img_array[29][18][7] <= img[13903];\
        in_img_array[29][18][8] <= img[13904];\
        in_img_array[29][18][9] <= img[13905];\
        in_img_array[29][18][10] <= img[13906];\
        in_img_array[29][18][11] <= img[13907];\
        in_img_array[29][18][12] <= img[13908];\
        in_img_array[29][18][13] <= img[13909];\
        in_img_array[29][18][14] <= img[13910];\
        in_img_array[29][18][15] <= img[13911];\
        in_img_array[29][18][16] <= img[13912];\
        in_img_array[29][18][17] <= img[13913];\
        in_img_array[29][19][0] <= img[13914];\
        in_img_array[29][19][1] <= img[13915];\
        in_img_array[29][19][2] <= img[13916];\
        in_img_array[29][19][3] <= img[13917];\
        in_img_array[29][19][4] <= img[13918];\
        in_img_array[29][19][5] <= img[13919];\
        in_img_array[29][19][6] <= img[13920];\
        in_img_array[29][19][7] <= img[13921];\
        in_img_array[29][19][8] <= img[13922];\
        in_img_array[29][19][9] <= img[13923];\
        in_img_array[29][19][10] <= img[13924];\
        in_img_array[29][19][11] <= img[13925];\
        in_img_array[29][19][12] <= img[13926];\
        in_img_array[29][19][13] <= img[13927];\
        in_img_array[29][19][14] <= img[13928];\
        in_img_array[29][19][15] <= img[13929];\
        in_img_array[29][19][16] <= img[13930];\
        in_img_array[29][19][17] <= img[13931];\
        in_img_array[29][20][0] <= img[13932];\
        in_img_array[29][20][1] <= img[13933];\
        in_img_array[29][20][2] <= img[13934];\
        in_img_array[29][20][3] <= img[13935];\
        in_img_array[29][20][4] <= img[13936];\
        in_img_array[29][20][5] <= img[13937];\
        in_img_array[29][20][6] <= img[13938];\
        in_img_array[29][20][7] <= img[13939];\
        in_img_array[29][20][8] <= img[13940];\
        in_img_array[29][20][9] <= img[13941];\
        in_img_array[29][20][10] <= img[13942];\
        in_img_array[29][20][11] <= img[13943];\
        in_img_array[29][20][12] <= img[13944];\
        in_img_array[29][20][13] <= img[13945];\
        in_img_array[29][20][14] <= img[13946];\
        in_img_array[29][20][15] <= img[13947];\
        in_img_array[29][20][16] <= img[13948];\
        in_img_array[29][20][17] <= img[13949];\
        in_img_array[29][21][0] <= img[13950];\
        in_img_array[29][21][1] <= img[13951];\
        in_img_array[29][21][2] <= img[13952];\
        in_img_array[29][21][3] <= img[13953];\
        in_img_array[29][21][4] <= img[13954];\
        in_img_array[29][21][5] <= img[13955];\
        in_img_array[29][21][6] <= img[13956];\
        in_img_array[29][21][7] <= img[13957];\
        in_img_array[29][21][8] <= img[13958];\
        in_img_array[29][21][9] <= img[13959];\
        in_img_array[29][21][10] <= img[13960];\
        in_img_array[29][21][11] <= img[13961];\
        in_img_array[29][21][12] <= img[13962];\
        in_img_array[29][21][13] <= img[13963];\
        in_img_array[29][21][14] <= img[13964];\
        in_img_array[29][21][15] <= img[13965];\
        in_img_array[29][21][16] <= img[13966];\
        in_img_array[29][21][17] <= img[13967];\
        in_img_array[29][22][0] <= img[13968];\
        in_img_array[29][22][1] <= img[13969];\
        in_img_array[29][22][2] <= img[13970];\
        in_img_array[29][22][3] <= img[13971];\
        in_img_array[29][22][4] <= img[13972];\
        in_img_array[29][22][5] <= img[13973];\
        in_img_array[29][22][6] <= img[13974];\
        in_img_array[29][22][7] <= img[13975];\
        in_img_array[29][22][8] <= img[13976];\
        in_img_array[29][22][9] <= img[13977];\
        in_img_array[29][22][10] <= img[13978];\
        in_img_array[29][22][11] <= img[13979];\
        in_img_array[29][22][12] <= img[13980];\
        in_img_array[29][22][13] <= img[13981];\
        in_img_array[29][22][14] <= img[13982];\
        in_img_array[29][22][15] <= img[13983];\
        in_img_array[29][22][16] <= img[13984];\
        in_img_array[29][22][17] <= img[13985];\
        in_img_array[29][23][0] <= img[13986];\
        in_img_array[29][23][1] <= img[13987];\
        in_img_array[29][23][2] <= img[13988];\
        in_img_array[29][23][3] <= img[13989];\
        in_img_array[29][23][4] <= img[13990];\
        in_img_array[29][23][5] <= img[13991];\
        in_img_array[29][23][6] <= img[13992];\
        in_img_array[29][23][7] <= img[13993];\
        in_img_array[29][23][8] <= img[13994];\
        in_img_array[29][23][9] <= img[13995];\
        in_img_array[29][23][10] <= img[13996];\
        in_img_array[29][23][11] <= img[13997];\
        in_img_array[29][23][12] <= img[13998];\
        in_img_array[29][23][13] <= img[13999];\
        in_img_array[29][23][14] <= img[14000];\
        in_img_array[29][23][15] <= img[14001];\
        in_img_array[29][23][16] <= img[14002];\
        in_img_array[29][23][17] <= img[14003];\
        in_img_array[29][24][0] <= img[14004];\
        in_img_array[29][24][1] <= img[14005];\
        in_img_array[29][24][2] <= img[14006];\
        in_img_array[29][24][3] <= img[14007];\
        in_img_array[29][24][4] <= img[14008];\
        in_img_array[29][24][5] <= img[14009];\
        in_img_array[29][24][6] <= img[14010];\
        in_img_array[29][24][7] <= img[14011];\
        in_img_array[29][24][8] <= img[14012];\
        in_img_array[29][24][9] <= img[14013];\
        in_img_array[29][24][10] <= img[14014];\
        in_img_array[29][24][11] <= img[14015];\
        in_img_array[29][24][12] <= img[14016];\
        in_img_array[29][24][13] <= img[14017];\
        in_img_array[29][24][14] <= img[14018];\
        in_img_array[29][24][15] <= img[14019];\
        in_img_array[29][24][16] <= img[14020];\
        in_img_array[29][24][17] <= img[14021];\
        in_img_array[29][25][0] <= img[14022];\
        in_img_array[29][25][1] <= img[14023];\
        in_img_array[29][25][2] <= img[14024];\
        in_img_array[29][25][3] <= img[14025];\
        in_img_array[29][25][4] <= img[14026];\
        in_img_array[29][25][5] <= img[14027];\
        in_img_array[29][25][6] <= img[14028];\
        in_img_array[29][25][7] <= img[14029];\
        in_img_array[29][25][8] <= img[14030];\
        in_img_array[29][25][9] <= img[14031];\
        in_img_array[29][25][10] <= img[14032];\
        in_img_array[29][25][11] <= img[14033];\
        in_img_array[29][25][12] <= img[14034];\
        in_img_array[29][25][13] <= img[14035];\
        in_img_array[29][25][14] <= img[14036];\
        in_img_array[29][25][15] <= img[14037];\
        in_img_array[29][25][16] <= img[14038];\
        in_img_array[29][25][17] <= img[14039];\
        in_img_array[29][26][0] <= img[14040];\
        in_img_array[29][26][1] <= img[14041];\
        in_img_array[29][26][2] <= img[14042];\
        in_img_array[29][26][3] <= img[14043];\
        in_img_array[29][26][4] <= img[14044];\
        in_img_array[29][26][5] <= img[14045];\
        in_img_array[29][26][6] <= img[14046];\
        in_img_array[29][26][7] <= img[14047];\
        in_img_array[29][26][8] <= img[14048];\
        in_img_array[29][26][9] <= img[14049];\
        in_img_array[29][26][10] <= img[14050];\
        in_img_array[29][26][11] <= img[14051];\
        in_img_array[29][26][12] <= img[14052];\
        in_img_array[29][26][13] <= img[14053];\
        in_img_array[29][26][14] <= img[14054];\
        in_img_array[29][26][15] <= img[14055];\
        in_img_array[29][26][16] <= img[14056];\
        in_img_array[29][26][17] <= img[14057];\
        in_img_array[29][27][0] <= img[14058];\
        in_img_array[29][27][1] <= img[14059];\
        in_img_array[29][27][2] <= img[14060];\
        in_img_array[29][27][3] <= img[14061];\
        in_img_array[29][27][4] <= img[14062];\
        in_img_array[29][27][5] <= img[14063];\
        in_img_array[29][27][6] <= img[14064];\
        in_img_array[29][27][7] <= img[14065];\
        in_img_array[29][27][8] <= img[14066];\
        in_img_array[29][27][9] <= img[14067];\
        in_img_array[29][27][10] <= img[14068];\
        in_img_array[29][27][11] <= img[14069];\
        in_img_array[29][27][12] <= img[14070];\
        in_img_array[29][27][13] <= img[14071];\
        in_img_array[29][27][14] <= img[14072];\
        in_img_array[29][27][15] <= img[14073];\
        in_img_array[29][27][16] <= img[14074];\
        in_img_array[29][27][17] <= img[14075];\
        in_img_array[29][28][0] <= img[14076];\
        in_img_array[29][28][1] <= img[14077];\
        in_img_array[29][28][2] <= img[14078];\
        in_img_array[29][28][3] <= img[14079];\
        in_img_array[29][28][4] <= img[14080];\
        in_img_array[29][28][5] <= img[14081];\
        in_img_array[29][28][6] <= img[14082];\
        in_img_array[29][28][7] <= img[14083];\
        in_img_array[29][28][8] <= img[14084];\
        in_img_array[29][28][9] <= img[14085];\
        in_img_array[29][28][10] <= img[14086];\
        in_img_array[29][28][11] <= img[14087];\
        in_img_array[29][28][12] <= img[14088];\
        in_img_array[29][28][13] <= img[14089];\
        in_img_array[29][28][14] <= img[14090];\
        in_img_array[29][28][15] <= img[14091];\
        in_img_array[29][28][16] <= img[14092];\
        in_img_array[29][28][17] <= img[14093];\
        in_img_array[29][29][0] <= img[14094];\
        in_img_array[29][29][1] <= img[14095];\
        in_img_array[29][29][2] <= img[14096];\
        in_img_array[29][29][3] <= img[14097];\
        in_img_array[29][29][4] <= img[14098];\
        in_img_array[29][29][5] <= img[14099];\
        in_img_array[29][29][6] <= img[14100];\
        in_img_array[29][29][7] <= img[14101];\
        in_img_array[29][29][8] <= img[14102];\
        in_img_array[29][29][9] <= img[14103];\
        in_img_array[29][29][10] <= img[14104];\
        in_img_array[29][29][11] <= img[14105];\
        in_img_array[29][29][12] <= img[14106];\
        in_img_array[29][29][13] <= img[14107];\
        in_img_array[29][29][14] <= img[14108];\
        in_img_array[29][29][15] <= img[14109];\
        in_img_array[29][29][16] <= img[14110];\
        in_img_array[29][29][17] <= img[14111];\
    end\
end